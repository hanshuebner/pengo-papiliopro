-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "747FB557CE90AA7D9D20080F7756C943A329C1212E6D756C94766C3D6F322F1D";
    attribute INIT_01 of inst : label is "E6DE95137F7BF7BEE4920E855FF0369DBB76ED818181010808090951A39DD1FF";
    attribute INIT_02 of inst : label is "DDF8C5DBD9BF8C7FA53657ED635B97F6BEB10FD0EEBD818BEB7E7CFA947E8007";
    attribute INIT_03 of inst : label is "F25AA23BEFA7FA8DBB6DA77F9CE3177FC99818726465F3030E4C0C3EFAF65ECB";
    attribute INIT_04 of inst : label is "D885B7225DB8F69877237180261C7B5D998038A0F64366CD9B37A183F26887E7";
    attribute INIT_05 of inst : label is "EDDB1D3ED51E27B31D15E8D7A35BA6E5EB96C2E6B2912BD9AEC33310B6216C42";
    attribute INIT_06 of inst : label is "6F61016CD9D3A474732FBED8FDB7D63755B3D90CE5308E90928402C6C6EFA2B6";
    attribute INIT_07 of inst : label is "76EDDBDBB76F6EDDBDBB76EABAA5114C13A510F64888F65BB76EDDBCDA6B18E3";
    attribute INIT_08 of inst : label is "ADCEDEC6BAE5D72F118E71ACCDF9C8A1CE3C99AC796E3CA11E58877287CFEDC6";
    attribute INIT_09 of inst : label is "8CC56A3AD9FA43A8F62073A660063FDA8B42B0DD65BC68237DFD9CC3C76777B2";
    attribute INIT_0A of inst : label is "3E945A1401D35877601C9D263FDA8B42B8F6D479A1D01A8BA548CD42B8ED9D12";
    attribute INIT_0B of inst : label is "0DC436F9F2EF5AD27C387A974C558BEE9757A17E5F8E7BDA6D369D361507BA8B";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFD55E2A2DDBB76EE21B7A0A9EF256F7C45C6C371B";
    attribute INIT_0D of inst : label is "2946294629462946294629462946294629462946294629462946294629462946";
    attribute INIT_0E of inst : label is "2946294629462946294629462946294629462946294629462946294629462946";
    attribute INIT_0F of inst : label is "2946294629462946294629462946294629462946294629462946294629462946";
    attribute INIT_10 of inst : label is "15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4";
    attribute INIT_11 of inst : label is "15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4";
    attribute INIT_12 of inst : label is "15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4";
    attribute INIT_13 of inst : label is "15B415B415B415B415B415B415B415B415B415B415B415B415B415B415B415B4";
    attribute INIT_14 of inst : label is "2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC";
    attribute INIT_15 of inst : label is "2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC";
    attribute INIT_16 of inst : label is "2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC";
    attribute INIT_17 of inst : label is "2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC2EEC";
    attribute INIT_18 of inst : label is "7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E";
    attribute INIT_19 of inst : label is "7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E";
    attribute INIT_1A of inst : label is "7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E";
    attribute INIT_1B of inst : label is "7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E7F2E";
    attribute INIT_1C of inst : label is "074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A";
    attribute INIT_1D of inst : label is "074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A";
    attribute INIT_1E of inst : label is "074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A";
    attribute INIT_1F of inst : label is "074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A074A";
    attribute INIT_20 of inst : label is "00081182008826000000110001080A000104080000800A000000000000000100";
    attribute INIT_21 of inst : label is "00C20ACF0000154F40A84A9C0088153301000A4F00980937818018D000802A3C";
    attribute INIT_22 of inst : label is "04080947040D0A9D05800D1B00400AB728220C2C001A295838300E70000809A3";
    attribute INIT_23 of inst : label is "07E1F84007E1F82000000A0201000C0006000A00040105000100002704010E0F";
    attribute INIT_24 of inst : label is "DE06DDBB400F3FFC000060BFFD03FFEE1CC03FFFFFFFFFFFFFFF185E15800000";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFBE000000000003FFFFC7401F7063803CDF";
    attribute INIT_26 of inst : label is "FFFFF1800000FF87FC80003FEFC4FFFC00003FFFFF7FF5FFFFFFFFDFF8000000";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAF80000000038001FFCF7FFFFFFF";
    attribute INIT_28 of inst : label is "FFB002100100901042108210810865BFFFEE836B772EFDFBFBF7FFF7FAFFFDFF";
    attribute INIT_29 of inst : label is "02AFBEFFFFFFFFF7FFFF556AA4914449529A291308445E56F7DEFDBAB52A4927";
    attribute INIT_2A of inst : label is "5555FEFFFFFFFFC00020000DFFFFFA6EFE2001C0049800000600001F54FFFF72";
    attribute INIT_2B of inst : label is "BDEFDEF78F7BDFBFBFBEFEFBEF7DEFDFEFF7FFBD9D2A949C924889042108410B";
    attribute INIT_2C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF9B";
    attribute INIT_2D of inst : label is "AAAAAAAA9010040200001008AFFF91BA13BB8ED0ACAB7636D2AD0A8AEEFDF7DF";
    attribute INIT_2E of inst : label is "FFFDFFEFFFFDFFF7BDAA0880495B7FBFFFFFFFFFFFFFFDF775EFEFEFBFFFFBFF";
    attribute INIT_2F of inst : label is "3AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA9FCFE";
    attribute INIT_30 of inst : label is "7E154327FFFFFFFFFFFFFFFDAAABFFFDAAAB6A0BFFF81A00FFFA1220FFF09220";
    attribute INIT_31 of inst : label is "C443903BFE50104BFFFFFF91111111111111111111111139FFFFFFF940401591";
    attribute INIT_32 of inst : label is "FFFFFFFF341041313041043331041031FFFFFFE0001BFF80049BFFFFFE111111";
    attribute INIT_33 of inst : label is "EC60606060726243FFFE44444449FFB0808080828080804BFFF8001BFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFF9100000E1FFFFFFF8411111E1FFFFFFFFAD5555E14C0000E30C0000E3";
    attribute INIT_35 of inst : label is "555005455154555555540155555005E1FFFFFFFFFFFFFFFFFFFFFFF8011111E1";
    attribute INIT_36 of inst : label is "5154555555540155555005E30014451555441515450511455541451555E10015";
    attribute INIT_37 of inst : label is "FFFFFFFFE0D54063E0D5406383050461FFFFFFFFFB3FEA41FFFF001555500545";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB054220D905040345157D4B1501540563";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC1515151551517440404040404040423";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC1504040540407551514040404040421";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFE4441093FFFFFFFFFFFFFFFFFFF9040410104091";
    attribute INIT_3E of inst : label is "6666666666CC150015001500150015E3FFFFFFFFFFFFFFFFFFFFFFFFFE400591";
    attribute INIT_3F of inst : label is "4400FFFFFFFFFFFF1504104104104161333333333315400550015000540015E1";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "11422FF95EA65D89264A2223590986655C4295757633909864A98950A2E35B71";
    attribute INIT_01 of inst : label is "8A0B2228014113C8018417088B45B9200000000C8C8C0C00000000050A004508";
    attribute INIT_02 of inst : label is "10F9133AB29FDA000FC598218A62D818C1C452C5898B352D8040BF7A695256B2";
    attribute INIT_03 of inst : label is "4503474013C9A336801004AAE739D7C51452D2A14B4A8A5A5429E9D3BC040180";
    attribute INIT_04 of inst : label is "011E080000E21A091001C40000710D048800E222B49B88102040893545219289";
    attribute INIT_05 of inst : label is "A34273CA6228D417A46623588D6093160C1830972666922BCD1A2823C047808F";
    attribute INIT_06 of inst : label is "40183F1512D819D158C4104BA69101A1980D6C72362138465C32E5989989CCD0";
    attribute INIT_07 of inst : label is "90A34242CD898A36262CD0AEDCDE03C60772890A13D080E08102040367B052B0";
    attribute INIT_08 of inst : label is "F1FF78EFC09800C376508A09DE1E664A11403BC07FBC3FDA1FED0BBF6207E434";
    attribute INIT_09 of inst : label is "15CE0442154D8A1110DAA2D8EDD46104D0642D10494157FEA4C2010A207FDE27";
    attribute INIT_0A of inst : label is "53668331696C12810DA916CE6144D0642D0808A6D504A4D0891AB6642D00C034";
    attribute INIT_0B of inst : label is "8011B800416318C464E9CC3891996CDA6E7A32EDE49CE044A6D12451972E0112";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFB880867102040808DC04BE25BF981410E4000000";
    attribute INIT_0D of inst : label is "44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0";
    attribute INIT_0E of inst : label is "44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0";
    attribute INIT_0F of inst : label is "44B044B044B044B044B044B044B044B044B044B044B044B044B044B044B044B0";
    attribute INIT_10 of inst : label is "89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF";
    attribute INIT_11 of inst : label is "89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF";
    attribute INIT_12 of inst : label is "89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF";
    attribute INIT_13 of inst : label is "89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF89AF";
    attribute INIT_14 of inst : label is "9425942594259425942594259425942594259425942594259425942594259425";
    attribute INIT_15 of inst : label is "9425942594259425942594259425942594259425942594259425942594259425";
    attribute INIT_16 of inst : label is "9425942594259425942594259425942594259425942594259425942594259425";
    attribute INIT_17 of inst : label is "9425942594259425942594259425942594259425942594259425942594259425";
    attribute INIT_18 of inst : label is "8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95";
    attribute INIT_19 of inst : label is "8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95";
    attribute INIT_1A of inst : label is "8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95";
    attribute INIT_1B of inst : label is "8A958A958A958A958A958A958A958A958A958A958A958A958A958A958A958A95";
    attribute INIT_1C of inst : label is "8233823382338233823382338233823382338233823382338233823382338233";
    attribute INIT_1D of inst : label is "8233823382338233823382338233823382338233823382338233823382338233";
    attribute INIT_1E of inst : label is "8233823382338233823382338233823382338233823382338233823382338233";
    attribute INIT_1F of inst : label is "8233823382338233823382338233823382338233823382338233823382338233";
    attribute INIT_20 of inst : label is "FF80037CFF0812FFFF8814FFFE8809FFFF800BFF7F040BFF0000000000000100";
    attribute INIT_21 of inst : label is "3F30134B7F90598F7F104D5D3EB007B47E1852507F1840477F0050C0FE002104";
    attribute INIT_22 of inst : label is "070825D907002013078006872342038F2782011C0FE006380FE825303FF83362";
    attribute INIT_23 of inst : label is "08E0E43C0071E01C00000BFC010009F002000DE0000006E2060101E4078103C0";
    attribute INIT_24 of inst : label is "DEF6C3293CCC87FA00007EB402BFFDE10245BFFFFFFFFFFFFD004541D5A0007F";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA40000000000040000193FE9001B909C1F";
    attribute INIT_26 of inst : label is "FFFFF003F8FE807C607BC23BE002100200003FE80079F1FFFFFFFFDFF800FFFF";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFA8400000401DA005FFF07FFFF7FF";
    attribute INIT_28 of inst : label is "001FFDFEFFFFFFFFFFFFFFFFEFFFBFFD30017EFFFFFFFFFFFFFFF7FFFFFFFFFF";
    attribute INIT_29 of inst : label is "F9504000002296BE7DEF7FFFFFFFFFFFFFFFFFFFEFFFF8FFFFFF7FFEDFFFFFFF";
    attribute INIT_2A of inst : label is "0000007F9B6DB6FFFFDFFFF3093FFBFFEFFFFFFFFFFFFFFFFFFFFFE300FFFFF7";
    attribute INIT_2B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEF3FFFF3FFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "000000000000000000000000000000000000000000000000000000000000003F";
    attribute INIT_2D of inst : label is "000000000FFFFFFFFFFFFFFFFBE463FFEC44712F5FFFFF3FFFF3FFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFE7FB6A48020AAF77FFFFFEFFFFFFFFFFFFFB7EEFF5B";
    attribute INIT_2F of inst : label is "550000000000000000000000000000000000000000000000000000000000003E";
    attribute INIT_30 of inst : label is "FFBBAC57FFFFFFFFFFFFFFFD2283FFFD0A234AA3FFFA92A0FFF89280FFF81280";
    attribute INIT_31 of inst : label is "AA1FC04DFF90109FFFFFFFD414141414141414141414140DFFFFFFFC2EAEAC6F";
    attribute INIT_32 of inst : label is "FFFFFFFF641041476041044561041045FFFFFFF4450DFFD1148DFFFFFF050505";
    attribute INIT_33 of inst : label is "F117711771155315FFFF0505051FFFC44CC44CC44CC44C1DFFFC088DFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFDEAAAAA1FFFFFFFFCFAEFFB1FFFFFFFFFBBFFFF17BAAAAA15BAAAAA17";
    attribute INIT_35 of inst : label is "451145511B16C50F9144516B45114597FFFFFFFFFFFFFFFFFFFFFFFCAAEFFB1F";
    attribute INIT_36 of inst : label is "1B16C50F9144516B45114597047F555145505B56D55FD554517F55514595047E";
    attribute INIT_37 of inst : label is "FFFFFFFFF0844095F0844095C24A0097FFFFFFFFFE91041FFFFF047E45114551";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEAFEDCE77E62EB9AAABD3A1B8AAE2AB9F";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFAAFFBDBBFBDAAABFEAAAAAAAAAA95";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFABFBBEEADAAEADAAABFEAAAAAAAAAA97";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFF9841065FFFFFFFFFFFFFFFFFFFD041410104067";
    attribute INIT_3E of inst : label is "6666666666CC405F555F550A000A0097FFFFFFFFFFFFFFFFFFFFFFFFFF800567";
    attribute INIT_3F of inst : label is "0100FFFFFFFFFFFF6836F3CF63A69A97333333333340404F4013D040A0102897";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "4933BAA95EF44F4DB52AAAAE0CCCEB69662655656C99CCCEB52CCDC89999EF78";
    attribute INIT_01 of inst : label is "1CDC733B2E1486E2418613882618BDB3972E5C880008000E060E0624C91924CE";
    attribute INIT_02 of inst : label is "C8D891A02A20171D8A66DDC9E9F35DFCEEF65390CFE5E4AE49EFFD78B324A527";
    attribute INIT_03 of inst : label is "AF6B6766FE5E1BBFE259228AA5294A2EBD4BCABD2F2AE97957A5E55C50BAD65A";
    attribute INIT_04 of inst : label is "C9CF96198C729F902318E50CC6394FC8118C72F7EDDBDE7CF9F2B887AF79171F";
    attribute INIT_05 of inst : label is "4C996CB7B33A1097B73779DDE779E7A74E9E50F7BFF0984BC9E91A39F273E4E7";
    attribute INIT_06 of inst : label is "6C2F0A6C18EB4DA3795C71C367D582B5FD17E56A5719B562C51626575665EAE7";
    attribute INIT_07 of inst : label is "074C991D326474C991D3267E8EEB102200E1019F587C12B9B366CD9EF7E95AF8";
    attribute INIT_08 of inst : label is "5C550009606C0763631CE885131F46639D10A262AFBD57DCABEE177F62000D59";
    attribute INIT_09 of inst : label is "BD9F0E6BC496C9399413B16EE9D27D96DB6BB5F77FE52A2229870519F32A8004";
    attribute INIT_0A of inst : label is "05B6DB5508B7DADD43258B6EFD96DB6BB5AF9CCB64B476DB7CDA5B6BBDBBFB15";
    attribute INIT_0B of inst : label is "BC95BE44715EF7BC01D7B02F19DDCE3EFD7FB4DFF17AD93FDB6DB3CD874D939B";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFBCD4ACFACD9B364ADF2F86B2F7DE5695F1E6F379";
    attribute INIT_0D of inst : label is "4000400040004000400040004000400040004000400040004000400040004000";
    attribute INIT_0E of inst : label is "4000400040004000400040004000400040004000400040004000400040004000";
    attribute INIT_0F of inst : label is "4000400040004000400040004000400040004000400040004000400040004000";
    attribute INIT_10 of inst : label is "0736073607360736073607360736073607360736073607360736073607360736";
    attribute INIT_11 of inst : label is "0736073607360736073607360736073607360736073607360736073607360736";
    attribute INIT_12 of inst : label is "0736073607360736073607360736073607360736073607360736073607360736";
    attribute INIT_13 of inst : label is "0736073607360736073607360736073607360736073607360736073607360736";
    attribute INIT_14 of inst : label is "34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA";
    attribute INIT_15 of inst : label is "34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA";
    attribute INIT_16 of inst : label is "34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA";
    attribute INIT_17 of inst : label is "34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA34FA";
    attribute INIT_18 of inst : label is "3080308030803080308030803080308030803080308030803080308030803080";
    attribute INIT_19 of inst : label is "3080308030803080308030803080308030803080308030803080308030803080";
    attribute INIT_1A of inst : label is "3080308030803080308030803080308030803080308030803080308030803080";
    attribute INIT_1B of inst : label is "3080308030803080308030803080308030803080308030803080308030803080";
    attribute INIT_1C of inst : label is "0310031003100310031003100310031003100310031003100310031003100310";
    attribute INIT_1D of inst : label is "0310031003100310031003100310031003100310031003100310031003100310";
    attribute INIT_1E of inst : label is "0310031003100310031003100310031003100310031003100310031003100310";
    attribute INIT_1F of inst : label is "0310031003100310031003100310031003100310031003100310031003100310";
    attribute INIT_20 of inst : label is "0008330200083600000814000008080081800800008008000000000000000100";
    attribute INIT_21 of inst : label is "0042120800005050000040E3410048C801804DA001804187819843FF00081303";
    attribute INIT_22 of inst : label is "040121680085206000882040200A2440206A268110280480102A0600000A3201";
    attribute INIT_23 of inst : label is "388003C0300007E000000C0501000E0F05000E1F0200073E0400013C04800278";
    attribute INIT_24 of inst : label is "0000004000001002000210000001000200008000000000000000000888000040";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000000000004080820000001000";
    attribute INIT_26 of inst : label is "0012000202025000400000000000000000000080000020000000000000004000";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0200000000080000010000000008";
    attribute INIT_28 of inst : label is "00104211010010104210A210910865FD10117F9488D102040408080805000203";
    attribute INIT_29 of inst : label is "FD524000002296BE7FFFD52AA493444952922913184559AD0821824555AA4927";
    attribute INIT_2A of inst : label is "000000004000003FFFDFFFE20937FE6EFE2001C00C980000060000030000008D";
    attribute INIT_2B of inst : label is "42102108608420404041010410821020100C00426DEA949C924889C42108410B";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000004";
    attribute INIT_2D of inst : label is "000000000010040200001008AFE46245EC44412F535489C92D5EF57511020823";
    attribute INIT_2E of inst : label is "00020010000200084255F7FFB6A48020AAF77FFFFFEFFDF775EFEDEFF7FEFF5B";
    attribute INIT_2F of inst : label is "0500000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "7E015077FFFFFFFFFFFFFFFD2003FFFD00234003FFF89A28FFF89A28FFF89A28";
    attribute INIT_31 of inst : label is "40159A4FFE54541FFFFFFF8015400015400015400015400DFFFFFFFBD0505645";
    attribute INIT_32 of inst : label is "FFFFFFFF1FBEFB4F1EFBEF4D1BEFBE4DFFFFFFE4E70FFF939C8FFFFFFE005500";
    attribute INIT_33 of inst : label is "E511177771333317FFFE0550021DFF94444CCCC6444CCC1DFFF8AA8FFFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFF95400009FFFFFFFF90114559FFFFFFFFF2555559D4555559D0400009F";
    attribute INIT_35 of inst : label is "AFAAAAABA0B82EADABEAAAA2AFAAAA1DFFFFFFFFFFFFFFFFFFFFFFF80114559F";
    attribute INIT_36 of inst : label is "A0B82EADABEAAAA2AFAAAA1D0277EABAAFEBE1FC6BBDFAAEABF7EABAAF1D0276";
    attribute INIT_37 of inst : label is "FFFFFFFFEA7CEA17EA7CEA17A9B7EA17FFFFFFFFF9015015FFFF0276AFAAAAAB";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFB1111555555C44541110000024449111D";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC404015155151544040551515151515D";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFEC515115155151544040440404040405F";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFE44EBF45FFFFFFFFFFFFFFFFFFF9EFA7BE9EFA45";
    attribute INIT_3E of inst : label is "6666666666CC3FA03FA03FA03FA03F15FFFFFFFFFFFFFFFFFFFFFFFFFE5AEF47";
    attribute INIT_3F of inst : label is "1401FFFFFFFFFFFF17CD1C718C18619733333333333FEEA5FBA97EAA5FAA9715";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "C7D19006F57FEA6671DD00039DFD61B299D7EA9A85E76666F2FF66BC61DAA5B0";
    attribute INIT_01 of inst : label is "348D888322BF01257AE9A9C0737303AA97363FAAD5D5AAA85657A8A2C7DFE2E2";
    attribute INIT_02 of inst : label is "5BADEB80EF0A09ACFFD967AEA4F5E7A6839B28FA5786838AE783575278F6BBA3";
    attribute INIT_03 of inst : label is "D2CEB1AB4B757BA83E793C08ED7BC2864BB5400BD4D42A8AABDA2A0E43F52191";
    attribute INIT_04 of inst : label is "CEFE87AAAAB4E2EA3AAA71C488946A60EAEE34A23DDF2E2EFADB27E978668BC5";
    attribute INIT_05 of inst : label is "BD7AA9A1B55BC44E5C4C910299484180A9530ABCF6BD1DFB86F7228C91950230";
    attribute INIT_06 of inst : label is "DC5B80FA07DBC0E1D30661A86DBCD6367B39B9C8FF5BCF839EB7AB271620BAAF";
    attribute INIT_07 of inst : label is "3EBD0686F56B99E2ADAF81BF7BB3AA21077F20AA3C9D86047375FA00FB699A97";
    attribute INIT_08 of inst : label is "F8EE8129F554DFF7FF0993CE8B07AAB6C8D3E6352DBA43864B6F522ED6D50A79";
    attribute INIT_09 of inst : label is "4F75EEF959F7BABBA52902E8F547238B0DD08EC0F8B4AAAA5AEDFAB2F2A23540";
    attribute INIT_0A of inst : label is "97576C8EFFDD6A66FAB6F9FF9E29A9B27A7EE679DB131BA9DDEBF9B27A61A98B";
    attribute INIT_0B of inst : label is "BC8F013BAEBD3603977F3ABF1F56466257D6D0A65FEF24AEFF75A820199F4BB8";
    attribute INIT_0C of inst : label is "0000555500005555000055557FCD3AAF47FD2E4389906936D9FF69C6F7EEBA39";
    attribute INIT_0D of inst : label is "54A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA02";
    attribute INIT_0E of inst : label is "7C0028007C0028007C0028007C0028007C0028007C0028007C0028007C002800";
    attribute INIT_0F of inst : label is "54A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA0254A8AA02";
    attribute INIT_10 of inst : label is "4AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B6";
    attribute INIT_11 of inst : label is "4AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E58";
    attribute INIT_12 of inst : label is "4AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B64AEB95B6";
    attribute INIT_13 of inst : label is "4AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E584AEB7E58";
    attribute INIT_14 of inst : label is "6BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB9674";
    attribute INIT_15 of inst : label is "6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E";
    attribute INIT_16 of inst : label is "6BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB96746BAB9674";
    attribute INIT_17 of inst : label is "6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E6BAB6D9E";
    attribute INIT_18 of inst : label is "2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C";
    attribute INIT_19 of inst : label is "2AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB5572";
    attribute INIT_1A of inst : label is "2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C2AEBFF9C";
    attribute INIT_1B of inst : label is "2AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB55722AEB5572";
    attribute INIT_1C of inst : label is "522B857C522B857C522B857C522B857C522B857C522B857C522B857C522B857C";
    attribute INIT_1D of inst : label is "522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82";
    attribute INIT_1E of inst : label is "522B857C522B857C522B857C522B857C522B857C522B857C522B857C522B857C";
    attribute INIT_1F of inst : label is "522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82522B7B82";
    attribute INIT_20 of inst : label is "FF77A829FF77A8AAFF77A8AAFF77A0AA7FF3A0AAFF7BA0AAFFFFAAAAFFFFABAA";
    attribute INIT_21 of inst : label is "551FA9EE157DABFA157DAA49157DAA66555DAA1A554DAA67554DAB7A55DDAAD6";
    attribute INIT_22 of inst : label is "FF73AAFBFFFFAAB8FF7FAAAEFFB7AAA2FF97AAF9DFC7ABEEDFC7ABAAFFE7ABF9";
    attribute INIT_23 of inst : label is "5DC48EEA5DC58E8A5555A2AC5555A2AA5555A2BA5555AA895555AA8E55D5AAEA";
    attribute INIT_24 of inst : label is "210D5FF561117951FFFFD5F7FEC2555FFFAD55550000555501FFFFFF162FAAD5";
    attribute INIT_25 of inst : label is "AAAA5555AAAA5555AAAA5555AAAA55145555AAAA55FF5555FBAA55547EFF5475";
    attribute INIT_26 of inst : label is "0000579F0785FFD78B4447D70FFAFFFDFFFFD55FFF8757550000557583DFD555";
    attribute INIT_27 of inst : label is "AAAA5555AAAA5555AAAA5555AAAA5555AAAA0555FFFB6AA5FFFC55552AAA5155";
    attribute INIT_28 of inst : label is "FFFFEAABFFFFAAAAFFFFAAAAFFFFEAEAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAA";
    attribute INIT_29 of inst : label is "5157AAAA5555AAA257552AEA5557BAAA555DAAA85555AAAE5555AAAB5555AAAB";
    attribute INIT_2A of inst : label is "FFFFABAABFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAABFFFFAAAA";
    attribute INIT_2B of inst : label is "5555AAAA7555AAAA5555AAAA5555AAAA5553AAAA5555AAAE5555AAEA5555AAAB";
    attribute INIT_2C of inst : label is "FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAEA";
    attribute INIT_2D of inst : label is "5555AAAA5555AAAA5555AAAA5555A2AA7555BAAA5555AAEA5555AABA5555AAAB";
    attribute INIT_2E of inst : label is "FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFABAAFFFFAAAB";
    attribute INIT_2F of inst : label is "0055AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAB";
    attribute INIT_30 of inst : label is "55FF00025555AAAA5555AAA84441AAA851010546555005745550443055504574";
    attribute INIT_31 of inst : label is "EAFF2FE255FFFFB25555002AFFFFEABFFFEABFFFAAAAFFE255550003FFFFFEE2";
    attribute INIT_32 of inst : label is "5555AAAAFFFF5500FFFE5500FFFA55005555AAA2FFFFAA88FEBFAAAA55AA5555";
    attribute INIT_33 of inst : label is "5FBBEEEEBBBB8CBA5555AFFFAAFF002BEEEEBBB3EEEE33B25556BEEA55550000";
    attribute INIT_34 of inst : label is "5555AAABAAEB51005555AAAAFEEB51005555AAAA1EFB5100FEFB5100FEFB5100";
    attribute INIT_35 of inst : label is "AAAFFABBAEABAEAFAAABFEAAAAAFFABA555500005555000055550001AAEBFFBA";
    attribute INIT_36 of inst : label is "AEAB5555AAAB0155AAAF0500AFEA5555AAAA5555AAAA5555AAAA5555AAFF5015";
    attribute INIT_37 of inst : label is "555500005FFFFFB25FFFFFB26BAAFBB25555000057FFFFB25555FAFEAAAFFABB";
    attribute INIT_38 of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAAFFFF0000FFFF0000FFFF1440FFFF0000";
    attribute INIT_39 of inst : label is "555500005555000055550000555500007FBFAFFFBFFBFFBFBBBBFBFBBBBBFBFA";
    attribute INIT_3A of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA7BBB4444BFBB4415AAAB4444BBBB4440";
    attribute INIT_3B of inst : label is "5555000055550000555500005555000055550000555500005555000055550000";
    attribute INIT_3C of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA";
    attribute INIT_3D of inst : label is "5555000055550000555500005FFBFFE255550000555500005557EFEFFFEBFFE2";
    attribute INIT_3E of inst : label is "CCCC3333CC661455AAAAD555AAAAD5085555AAAA5555AAAA5555AAAA55FF0508";
    attribute INIT_3F of inst : label is "FEAB000055550000EBAAFFFFAAAAFFB29999CCCC99EBEEEFAEEEFEEEAAEEBFB2";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "B9B8FA8450310E01064088882CCCCB446608413130D9CCCCB08CC80E1C116C08";
    attribute INIT_01 of inst : label is "2D41B77C2B60B8E4575F73BA80649C90102040848484040606060602855AE6E2";
    attribute INIT_02 of inst : label is "30D6182522A0121548081D51C5741D5CEAE777A610F1E2E69B6AC08524A135E0";
    attribute INIT_03 of inst : label is "1790646C58AC81DB601001FC11846A805E2BAB80AEAE05757015D5C0104DC9B9";
    attribute INIT_04 of inst : label is "898F18BB99CF1DB367339E5DCCE78ED9B399CF0006E9C0408102181417BD702C";
    attribute INIT_05 of inst : label is "12246A03C3305B547777FB9FEE71FCE7CFDC5301C3A2BD8AABA50C31E263C4C7";
    attribute INIT_06 of inst : label is "404A0410810451A082504903500B64A0A624321307013543721B91018191E4E9";
    attribute INIT_07 of inst : label is "0912242408101120404089104EECF6FDFD8C6400514514C142850A1427D26124";
    attribute INIT_08 of inst : label is "53772B1D4C82641072DEF941128F0C5BDF2922532C459620CB10699884371522";
    attribute INIT_09 of inst : label is "58AA066848824919C25380260A934D961B45B5D385C12022861B6CA902BB8ACD";
    attribute INIT_0A of inst : label is "6090DA233812DACC250781214D961B45B58D8CC130A4121B0A304905B59ADB00";
    attribute INIT_0B of inst : label is "509A9C59155294A48250A64009DC6E5CF51F825EF04AD10B45A2D041242D1198";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF9CCBC4780810204D4E2014A8CFDC557AF68742A1";
    attribute INIT_0D of inst : label is "11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE";
    attribute INIT_0E of inst : label is "11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE";
    attribute INIT_0F of inst : label is "11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE11FE";
    attribute INIT_10 of inst : label is "8811881188118811881188118811881188118811881188118811881188118811";
    attribute INIT_11 of inst : label is "8811881188118811881188118811881188118811881188118811881188118811";
    attribute INIT_12 of inst : label is "8811881188118811881188118811881188118811881188118811881188118811";
    attribute INIT_13 of inst : label is "8811881188118811881188118811881188118811881188118811881188118811";
    attribute INIT_14 of inst : label is "849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F";
    attribute INIT_15 of inst : label is "849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F";
    attribute INIT_16 of inst : label is "849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F";
    attribute INIT_17 of inst : label is "849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F849F";
    attribute INIT_18 of inst : label is "9011901190119011901190119011901190119011901190119011901190119011";
    attribute INIT_19 of inst : label is "9011901190119011901190119011901190119011901190119011901190119011";
    attribute INIT_1A of inst : label is "9011901190119011901190119011901190119011901190119011901190119011";
    attribute INIT_1B of inst : label is "9011901190119011901190119011901190119011901190119011901190119011";
    attribute INIT_1C of inst : label is "8003800380038003800380038003800380038003800380038003800380038003";
    attribute INIT_1D of inst : label is "8003800380038003800380038003800380038003800380038003800380038003";
    attribute INIT_1E of inst : label is "8003800380038003800380038003800380038003800380038003800380038003";
    attribute INIT_1F of inst : label is "8003800380038003800380038003800380038003800380038003800380038003";
    attribute INIT_20 of inst : label is "0000600300086500000005000100080000080900010008000000000000000000";
    attribute INIT_21 of inst : label is "00422240002044C0002044C3002004880000042000100087001000E001006040";
    attribute INIT_22 of inst : label is "0401060104050282048A06A4244206A8286206D318302560182227A0001207C3";
    attribute INIT_23 of inst : label is "001104000000000000000A0600000A0006010A00020102000401040404812600";
    attribute INIT_24 of inst : label is "DF03FD9BE00F5BF80000705DFEC3FFF61E503FFFFFFFFFFFFF7F585F0BC00000";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAE000000000001FFFFC3801F70F100AC7F";
    attribute INIT_26 of inst : label is "FFFFF98000047FC5F800083DF7E6F7FC00003FFFFF7EFFFFFFFFFFDF7C200000";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFAFC0000400038003FFCFFFFFFBFF";
    attribute INIT_28 of inst : label is "0008000000000000000020000000010020100100001000000000000000000001";
    attribute INIT_29 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2D of inst : label is "0000000010000000000000000400100020002000080000800008002000000002";
    attribute INIT_2E of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_2F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_30 of inst : label is "FF400157FFFFFFFFFFFFFFFFAEABFFFFBAABEEFBFFFABAAAFFFAFAAAFFFABAAA";
    attribute INIT_31 of inst : label is "5555F455FF400055FFFFFFD5555540000015555540000015FFFFFFFD00000055";
    attribute INIT_32 of inst : label is "FFFFFFFF554054555501505554054055FFFFFFF44555FFD55515FFFFFF000000";
    attribute INIT_33 of inst : label is "F511111111111555FFFF55555055FFD44444444444444455FFFC4555FFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFD54410455FFFFFFFC01145155FFFFFFFF350451555504515555045155";
    attribute INIT_35 of inst : label is "55500555515455555554015555500555FFFFFFFFFFFFFFFFFFFFFFFC01145155";
    attribute INIT_36 of inst : label is "5154555555540155555005550555505555555555515554155555505555550555";
    attribute INIT_37 of inst : label is "FFFFFFFFF5400455F5400455D5555555FFFFFFFFFD400055FFFF055555500555";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF50155555551155555555411455515555";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0404040540405444444444444444455";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD4040404144041511110000000000015";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFF7651555FFFFFFFFFFFFFFFFFFFF555840355555";
    attribute INIT_3E of inst : label is "6666666666CC41554055405540554055FFFFFFFFFFFFFFFFFFFFFFFFFF610555";
    attribute INIT_3F of inst : label is "5501FFFFFFFFFFFF410000000000005533333333334111100444011100444055";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "B52ED2AC54C53AF5EE37F7F2131355D7FE39D1216BF975754B3174FF3EE476E5";
    attribute INIT_01 of inst : label is "3971F77141DFE31AB1C7645FFC255C776051D455575755545555557D543C3D45";
    attribute INIT_02 of inst : label is "9C59C8C058555F2C822B954D164E1557EBF15D77B9F9939B9C6B682CE3B9C593";
    attribute INIT_03 of inst : label is "5590151514B984574D345001D4B57FF55601959806077D4D1DB03500548DCEC5";
    attribute INIT_04 of inst : label is "9FDCDBDD0067F69591FFFBD55DEDF97537443AFF653B7E5CEC66F447D7B85B37";
    attribute INIT_05 of inst : label is "8342155C46680AA16664C47755C61C1D9171C3C46567C2EF996CF1714D5DFDC4";
    attribute INIT_06 of inst : label is "FAB4D4452F7E0C78B4EDB2E79658EF5B9CC6E02B94C6BE56214EF2FE3A22273E";
    attribute INIT_07 of inst : label is "D0837B7B0D09ED6724209EC0141C85D4F4555847E17754BF0D1847F4678417E9";
    attribute INIT_08 of inst : label is "595582346FB1AE2566645497646CDD616546806457F0C01C55FD3CC0541D01A3";
    attribute INIT_09 of inst : label is "149E91131C65C54410559F1C1F703C61164D743F1D4F5FD5F51E3DD564FF8BBE";
    attribute INIT_0A of inst : label is "59CF4A87D1C74D762759477A51D61DD4C191D54F74E7529DB515DFD4C99E4DD2";
    attribute INIT_0B of inst : label is "D1795FDCCD47E4F0E441502D5198B15CEC595BD166505F7186517514656CB443";
    attribute INIT_0C of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAA9139A57F9CCA374A2E6FCF3B1F127BEFCDB3F279";
    attribute INIT_0D of inst : label is "D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400";
    attribute INIT_0E of inst : label is "55FD54A855FD54A855FD54A855FD54A855FD54A855FD54A855FD54A855FD54A8";
    attribute INIT_0F of inst : label is "D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400D7FF5400";
    attribute INIT_10 of inst : label is "AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555";
    attribute INIT_11 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_12 of inst : label is "AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555AAAAF555";
    attribute INIT_13 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_14 of inst : label is "AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555";
    attribute INIT_15 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_16 of inst : label is "AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555";
    attribute INIT_17 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_18 of inst : label is "AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555";
    attribute INIT_19 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_1A of inst : label is "AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555AAAAD555";
    attribute INIT_1B of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_1C of inst : label is "AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5";
    attribute INIT_1D of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_1E of inst : label is "AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5AAAAFDD5";
    attribute INIT_1F of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_20 of inst : label is "54DD555654DD515554DD535554DD5F5554555F5554555F555555555555555455";
    attribute INIT_21 of inst : label is "555D547D157D50D5157D51F6147D51DD545D51F554DD55DAD45D54F554DD55FD";
    attribute INIT_22 of inst : label is "50D5735454D577D754DD73D1715773DD7D5773C44D5551554D57535555577356";
    attribute INIT_23 of inst : label is "5DC471155DC57175555551535455515D51555155545551765055517150D5515D";
    attribute INIT_24 of inst : label is "8AAA9FAF2AAABEAFAAAA2BAFAAAAABAE8AABAAAAAAAAAAAAAAAA7A9FA8A5552A";
    attribute INIT_25 of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAA4B555555555500FFFF38AABEFF8C10BB6A";
    attribute INIT_26 of inst : label is "AAAAA6FEAAAABFAFAAEA9FEAAA9AFFFEAAAAEABFAA2BA4AAAAAAAA8AAA9AAAAA";
    attribute INIT_27 of inst : label is "AAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA57FF0000955AB008AAAF2AAAAEAA";
    attribute INIT_28 of inst : label is "550557555555D55551557555455555555555575555D5555555555D5551555557";
    attribute INIT_29 of inst : label is "555555555555555D5555D5555555555555555555455455555555555555555555";
    attribute INIT_2A of inst : label is "555555555555555555555555555555555555555555555555555555555555555D";
    attribute INIT_2B of inst : label is "5555555565555555555555555555555555555555551555555555555555555555";
    attribute INIT_2C of inst : label is "5555555555555555555555555555555555555555555555555555555555555555";
    attribute INIT_2D of inst : label is "5555555555555555555555555555555545555555515555555551555555555555";
    attribute INIT_2E of inst : label is "5555555555555555555554D55555557555555555555D555515555555755D5755";
    attribute INIT_2F of inst : label is "0155555555555555555555555555555555555555555555555555555555555755";
    attribute INIT_30 of inst : label is "55AA54025555AAAA5555AAAAEFA9AAAAFEA9ABFA555EAEBE555AEAAE555EAABE";
    attribute INIT_31 of inst : label is "EAFF2FAA55EAFFAA5555003FAAAAFFFFAAAAFFFFAAAAFFEA55550003AAAAFFAA";
    attribute INIT_32 of inst : label is "5555AAAAFAAA5500FAAA5500FAAA55005555AAA1EFBFAA84BEBFAAAA55AA5555";
    attribute INIT_33 of inst : label is "5FBBEEEEBBBBEEAA5555FFFFAAFF002BEEEEBBBBEEEEBBAA5556BEEA55550000";
    attribute INIT_34 of inst : label is "5555AAA9AAEB51005555AAA9AAAA55005555AAAA9EAA5500BEAA5500BEAA5500";
    attribute INIT_35 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFAA555500005555000055550003AAAAFFAA";
    attribute INIT_36 of inst : label is "AAAA5555AAAA5555AAAA5500AFEA5555AAAA5555AAAA5555AAAA5555AAFF5015";
    attribute INIT_37 of inst : label is "555500005AEAFFAA5AEAFFAA6BAAFFAA5555000057AAFFAA5555FABFAAAAFFFF";
    attribute INIT_38 of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAAEAAA5555AFAA5405AAAA5555AAAA5540";
    attribute INIT_39 of inst : label is "555500005555000055550000555500007AAAFFFFBEAAFEBFAAAAFFFFAAAAFFEA";
    attribute INIT_3A of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA7AAA5555BEAA5415AAAA5555AAAA5540";
    attribute INIT_3B of inst : label is "5555000055550000555500005555000055550000555500005555000055550000";
    attribute INIT_3C of inst : label is "5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA5555AAAA";
    attribute INIT_3D of inst : label is "5555000055550000555500005FEBFFAA55550000555500005556EFEFEAABFFAA";
    attribute INIT_3E of inst : label is "CCCC3333CC661455AAAA5555AAAA55005555AAAA5555AAAA5555AAAA55EB5500";
    attribute INIT_3F of inst : label is "AEAB000055550000EBAAFFFFAAAAFFAA9999CCCC99EBEEEFAEEEFEEEAAEEBFAA";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "717BBAAA403022FEFBFF77718E46C3A223BEFEDED39C646C384476DC49B16C20";
    attribute INIT_01 of inst : label is "8FC631163EB769786AA2A8C55182CDBD5AB4688000000000000000458BC5C5EF";
    attribute INIT_02 of inst : label is "9F54EF85098018A41FF247FC4B1907C63E200BCBE425C5C3DB7EE1C7FF77D6E1";
    attribute INIT_03 of inst : label is "C6ED7577D94FB8CB32492601BDEF75531B9C5C327170D38B864E2E1BEB2664CC";
    attribute INIT_04 of inst : label is "888B1388449DC4C180013BC4224EE260C0009DF59CECFD7AF1E32180C6CD398C";
    attribute INIT_05 of inst : label is "F9F3DFFCB1120A10B919488522112DA1428440C990B00D28CDDB37116A22D445";
    attribute INIT_06 of inst : label is "BF6300F848EF416A631C79C2F1C4D65FCBB0C79841F2EE03661B30F4F4CF3A3C";
    attribute INIT_07 of inst : label is "BCF9F3F3E7CFCF9F3F3E7CEBE323007001F008E60809F631AB568D1DF24B98EB";
    attribute INIT_08 of inst : label is "5D77AE057BE0DF053221081E222984442103C4462AC115608AB14DD580680C44";
    attribute INIT_09 of inst : label is "9D46A239C5D6CB88E600336F809625C759A0B59161D17F75FA63D45B8B3BAB81";
    attribute INIT_0A of inst : label is "15BACD0401B65AE6602C9B68258759A0B5C4C46B65903759E1C2DBA0B5C91B11";
    attribute INIT_0B of inst : label is "28EECC7078FBDEF31FBF606E9C4603AC33ACD1B6BFF7B5F6FB7DBD343B1B1889";
    attribute INIT_0C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFC467745EAD5A347766320312C24468EEB954AA51";
    attribute INIT_0D of inst : label is "7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00";
    attribute INIT_0E of inst : label is "7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00";
    attribute INIT_0F of inst : label is "7C007C007C007C007C007C007C007C007C007C007C007C007C007C007C007C00";
    attribute INIT_10 of inst : label is "1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE";
    attribute INIT_11 of inst : label is "1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE";
    attribute INIT_12 of inst : label is "1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE";
    attribute INIT_13 of inst : label is "1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE1FBE";
    attribute INIT_14 of inst : label is "3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE";
    attribute INIT_15 of inst : label is "3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE";
    attribute INIT_16 of inst : label is "3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE";
    attribute INIT_17 of inst : label is "3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE3EFE";
    attribute INIT_18 of inst : label is "7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE";
    attribute INIT_19 of inst : label is "7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE";
    attribute INIT_1A of inst : label is "7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE";
    attribute INIT_1B of inst : label is "7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE7FBE";
    attribute INIT_1C of inst : label is "077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E";
    attribute INIT_1D of inst : label is "077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E";
    attribute INIT_1E of inst : label is "077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E";
    attribute INIT_1F of inst : label is "077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E077E";
    attribute INIT_20 of inst : label is "00887880008078000088180000880000000C0000008400000000000000000000";
    attribute INIT_21 of inst : label is "004A396C002859D0002858E0002858C40008589000984848001859F0008878FC";
    attribute INIT_22 of inst : label is "008D2858008D2890008A28A0004A28A0006A28C0003A2964003A29A8001A39D0";
    attribute INIT_23 of inst : label is "0000000000000000000000000000000801010010040108200001082000812848";
    attribute INIT_24 of inst : label is "0000040040200100400000000000000002201000000000000000400010200000";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000000000008000000001000000000000";
    attribute INIT_26 of inst : label is "0000010000100020020004000008000000000000000401000000000042000000";
    attribute INIT_27 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0000002000000000002400003000";
    attribute INIT_28 of inst : label is "0048000000000000000020000000010020100100001000000000000000000001";
    attribute INIT_29 of inst : label is "0400010000000000801000000002000000000002000001000000800000800002";
    attribute INIT_2A of inst : label is "0000018040000000002000100008040010000000080000000000000281000000";
    attribute INIT_2B of inst : label is "0000000020000000000000000000000000040000008000080000008000000002";
    attribute INIT_2C of inst : label is "0000000000000000000000000000000000000000000000000000000000000060";
    attribute INIT_2D of inst : label is "0000000030000000000000000400100020002000080000800008002000000002";
    attribute INIT_2E of inst : label is "0000000000000000000001000000004000000000001000008000020040100402";
    attribute INIT_2F of inst : label is "D100000000000000000000000000000000000000000000000000000000020301";
    attribute INIT_30 of inst : label is "FF000157FFFFFFFFFFFFFFFFFFBBFFFFFEFBFBEFFFFABBEFFFFABEABFFFABAAB";
    attribute INIT_31 of inst : label is "4055D055FF400055FFFFFFC0000000000000000000000015FFFFFFFC00000055";
    attribute INIT_32 of inst : label is "FFFFFFFF500000555000005550000055FFFFFFF44515FFD11415FFFFFF000000";
    attribute INIT_33 of inst : label is "F511111111111155FFFF55555555FFD44444444444444455FFFD5115FFFFFFFF";
    attribute INIT_34 of inst : label is "FFFFFFFC00410455FFFFFFFC00000055FFFFFFFF340000551400005514000055";
    attribute INIT_35 of inst : label is "00000000000000000000000000000055FFFFFFFFFFFFFFFFFFFFFFFC00000055";
    attribute INIT_36 of inst : label is "0000000000000000000000550540000000000000000000000000000000550540";
    attribute INIT_37 of inst : label is "FFFFFFFFF0400055F0400055C1000055FFFFFFFFFD000055FFFF054000000000";
    attribute INIT_38 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF40000000050001500000144000000015";
    attribute INIT_39 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0000000140001400000000000000015";
    attribute INIT_3A of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFD0000000140001400000000000000015";
    attribute INIT_3B of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3C of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_3D of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFF5410055FFFFFFFFFFFFFFFFFFFC101040010055";
    attribute INIT_3E of inst : label is "6666666666CC55555555555555555555FFFFFFFFFFFFFFFFFFFFFFFFFF410055";
    attribute INIT_3F of inst : label is "4401FFFFFFFFFFFF410000000000005533333333334111100444011100444055";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "E0CFE5F7EA9BDC9A15827770B5FDB0AC898F2AAAFEB78A8B587F9A61E51BDBE7";
    attribute INIT_01 of inst : label is "0D9D611AAA02D07177D77DBFAE5C88EC932E19D70000575500005518D3C17489";
    attribute INIT_02 of inst : label is "57A31A7FEB2A96537D8CAAA2FDF5EAA9809432275696565D63801E7E3EC74340";
    attribute INIT_03 of inst : label is "A748656F5E0C5D9E335DE2009CC6354B9D9FCAAB7E7FABDBD67F6F69437F61DA";
    attribute INIT_04 of inst : label is "6235685511532B1DC5DD9A0055778CA41D550655CE6719A333D9C33E0DE5E0F2";
    attribute INIT_05 of inst : label is "DFFB0C39B11754407D57DDCF227964BBD7BE540DF0F9DD9C1DA75A157227D455";
    attribute INIT_06 of inst : label is "9A8766B2B2CEFC978DE0DF5F7FF62D234CDF58E46BFE30F6C8E9FD194C45CDC1";
    attribute INIT_07 of inst : label is "3EDF87873FEF1CA8BFB3A1C4226BFCD500404A09DC528FC432E4BC42B65F5821";
    attribute INIT_08 of inst : label is "BDBF79F7F36C28D841745762B9133B9175B219D97AE6FE8F0AB8FBBA68CAE6B7";
    attribute INIT_09 of inst : label is "9CDB777A45B2BEDDB517A5391AA651F61954C5C420E628285193C92E1B8AF58D";
    attribute INIT_0A of inst : label is "A61E3249263CB318FBE7B6DAEE5CB6AF3B6E3BA48F7CCCB6917E36AF3B67F67F";
    attribute INIT_0B of inst : label is "5CD4893C6D9D12070672255C8D767621FF5C96A67D67A483C97CEA6954B34DDA";
    attribute INIT_0C of inst : label is "5555000055550000555500007FF48BB36539C198CD193E09EDFC966B51CF8D26";
    attribute INIT_0D of inst : label is "444493BB444493BB444493BB444493BB444493BB444493BB444493BB444493BB";
    attribute INIT_0E of inst : label is "EEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBBEEEEBBBB";
    attribute INIT_0F of inst : label is "444493BB444493BB444493BB444493BB444493BB444493BB444493BB444493BB";
    attribute INIT_10 of inst : label is "D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105";
    attribute INIT_11 of inst : label is "D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041";
    attribute INIT_12 of inst : label is "D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105D4F20105";
    attribute INIT_13 of inst : label is "D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041D4F2E041";
    attribute INIT_14 of inst : label is "C7341041C7341041C7341041C7341041C7341041C7341041C7341041C7341041";
    attribute INIT_15 of inst : label is "C734C101C734C101C734C101C734C101C734C101C734C101C734C101C734C101";
    attribute INIT_16 of inst : label is "C7341041C7341041C7341041C7341041C7341041C7341041C7341041C7341041";
    attribute INIT_17 of inst : label is "C734C101C734C101C734C101C734C101C734C101C734C101C734C101C734C101";
    attribute INIT_18 of inst : label is "FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005";
    attribute INIT_19 of inst : label is "FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041";
    attribute INIT_1A of inst : label is "FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005FFD80005";
    attribute INIT_1B of inst : label is "FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041FFD88041";
    attribute INIT_1C of inst : label is "D1280455D1280455D1280455D1280455D1280455D1280455D1280455D1280455";
    attribute INIT_1D of inst : label is "D128F881D128F881D128F881D128F881D128F881D128F881D128F881D128F881";
    attribute INIT_1E of inst : label is "D1280455D1280455D1280455D1280455D1280455D1280455D1280455D1280455";
    attribute INIT_1F of inst : label is "D128F881D128F881D128F881D128F881D128F881D128F881D128F881D128F881";
    attribute INIT_20 of inst : label is "ABAAEE7CABAAEBFFABAAEBFFAAAAFFFF2B2AFFFFAA2AFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_21 of inst : label is "00C0555500805345000042570180021D01800275018014D78180074500004685";
    attribute INIT_22 of inst : label is "ABABFFA7ABAFFE6DABAAFE5B8E6AFF5782EAFF6D92AAFEDF92BAFE57AAAAFA7D";
    attribute INIT_23 of inst : label is "0880751508907175000059530000595503015955030151560101555101015515";
    attribute INIT_24 of inst : label is "545C0200544560005555002255150000F4D500005555000055D58000554AFF80";
    attribute INIT_25 of inst : label is "FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAE10000555500FD0000FFFFA801F97FC90A";
    attribute INIT_26 of inst : label is "5555004055D50002555500424D540801D555400055D500005555000051550000";
    attribute INIT_27 of inst : label is "FFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFF800FFFB1548EFEFAA00FFFFA2AA";
    attribute INIT_28 of inst : label is "AABABDFEAAAA7FFFAEAAFFFFBAAABEBFAAAAFDFFAA2AFFFFAAAAF7FFAEAAFFFD";
    attribute INIT_29 of inst : label is "0402555500005555021055150000455500085555100155510000555400005554";
    attribute INIT_2A of inst : label is "AAAAFFFFEAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFE2AAAFFF7";
    attribute INIT_2B of inst : label is "0000555510005555000055550000555500065555004055510000551500005554";
    attribute INIT_2C of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_2D of inst : label is "0000555520005555000055550600515510004555040055150004554500005554";
    attribute INIT_2E of inst : label is "AAAAFFFFAAAAFFFFAAAAFE7FAAAAFFDFAAAAFFFFAAA2FFFFEAAAFEFF8AA2FDFE";
    attribute INIT_2F of inst : label is "D000555500005555000055550000555500005555000055550000555500025555";
    attribute INIT_30 of inst : label is "AA410117AAAAFFFFAAAAFFFD5556FFFD55564003AAAF1000AAAF1000AAAF1000";
    attribute INIT_31 of inst : label is "1518F455AA155555AAAAFFD5155555555540000040150015AAAAFFFD55555555";
    attribute INIT_32 of inst : label is "AAAAFFFF055500150555001505550015AAAAFFF418C8FFD163C8FFFFAA550055";
    attribute INIT_33 of inst : label is "A044111142021155AAAA00005018FFD41111444499994455AAAB4115AAAAFFFF";
    attribute INIT_34 of inst : label is "AAAAFFFC55140445AAAAFFFC55550045AAAAFFFF615500454155004541550045";
    attribute INIT_35 of inst : label is "05055000041100000141540005055055AAAAFFFFAAAAFFFFAAAAFFFC55550455";
    attribute INIT_36 of inst : label is "0411515001410155050505455055050505551401515501410155050505100501";
    attribute INIT_37 of inst : label is "AAAAFFFFA5165555A516555594550055AAAAFFFFA8415555AAAA054005055000";
    attribute INIT_38 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFE11150000545500545100411554410445";
    attribute INIT_39 of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFC4041515515551515555111151511115";
    attribute INIT_3A of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFC5154000515500514445040451510405";
    attribute INIT_3B of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_3C of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFFAAAAFFFF";
    attribute INIT_3D of inst : label is "AAAAFFFFAAAAFFFFAAAAFFFFA2144055AAAAFFFFAAAAFFFFAAA9555515540055";
    attribute INIT_3E of inst : label is "3333666633994100D5550000D5550045AAAAFFFFAAAAFFFFAAAAFFFFAA140015";
    attribute INIT_3F of inst : label is "5054FFFFAAAAFFFF145500005555005566663333661411105111011155114055";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
