-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity ROM_PGM_0 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of ROM_PGM_0 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "5C2FDAAE2EDA2B3198CE6733102490476B6488DCA50900623E0000F6F948282D";
    attribute INIT_01 of inst : label is "0D1D6BB5DA6DBDF17DD0B2B0B0AE2BBA71C53548570BFF88D5238347948E24D6";
    attribute INIT_02 of inst : label is "7C6822100004650C4200008788408004518574C2B1C94C5E1FC5DC762ACD18B4";
    attribute INIT_03 of inst : label is "81809048681B99506A24674D074B6630B7BE5EAEEF663FF5F7DFFA71654FCFB9";
    attribute INIT_04 of inst : label is "4001709A0400B2B2C2F4857B380818DF28147D20A023228A014316947EA36404";
    attribute INIT_05 of inst : label is "0E423947A3D1E8E0B83CB8FB6AD6ED43F7EDE28B48845B6D92F6DEC19BDD056D";
    attribute INIT_06 of inst : label is "40E40285DC4B6F6862D1B6DFFBBFFE5FC2589992EC3D54D4ABBD8E8A04114DEA";
    attribute INIT_07 of inst : label is "EFB97C683DD1E0C90F04D8437EAAE8EA8DFF9F03252B53B59AC513D4CC890401";
    attribute INIT_08 of inst : label is "D37B8012926245C2932C0404A07210803115E8CA7DBE82369E88010B9BC88953";
    attribute INIT_09 of inst : label is "B6BB3412FDD043170C773EDDD20F5BF4957B3DCD31F34000046A75BEFDFB1377";
    attribute INIT_0A of inst : label is "0D20804820160EB48318AB23002B332DBEDBEDBEDADFAA70011761EC1C76DF7D";
    attribute INIT_0B of inst : label is "1F807917AD2051110868B22089064409A2C880241910268323830E7AE7A6C7B8";
    attribute INIT_0C of inst : label is "011729EF0ED6CE2A836715513A0812B1B6839990137AEA1909F682F5F390E600";
    attribute INIT_0D of inst : label is "8DB1B636C6D9FEF2F2F2AAAAA7A23F9F33C75EF6836C6D190A496C52B187AA70";
    attribute INIT_0E of inst : label is "65F7D8F6B3CDA0DE39C9E169364E8DDA5061A5F61B6F74F1A5249EFE7CE907EA";
    attribute INIT_0F of inst : label is "6638A714669BFDECA269BBFB28DACBEDB1D4F61C71C70CCD3D42B4A914090A4F";
    attribute INIT_10 of inst : label is "863FB76FB365196649CB724E1B8430E1A1B76C9ADF84E1276165F65B75BE4047";
    attribute INIT_11 of inst : label is "B42D03669B78C74BEB824EB8349C5759C534D142F15DC1A4E2BA29A2BAE97E2C";
    attribute INIT_12 of inst : label is "64FB7ED50E0E950E2E82901691499CBD2315492294EE4C1C11111AE41555777B";
    attribute INIT_13 of inst : label is "7788ED64A30CC1386E08C3304E1B8710DC219C8C71748DF43768A5DE36B9C932";
    attribute INIT_14 of inst : label is "9607AC6B009EC034600D883620C8A412090C82F2EED115AE9DE23B593B4456B2";
    attribute INIT_15 of inst : label is "3346E8CC69EC6DB4DC1B766E9BD775A205229F70453FDA408836BA5FE03BA769";
    attribute INIT_16 of inst : label is "E0D44B53A1C20CB8D74BD03F55D140861440068CE10180C0203004A2834CD1BA";
    attribute INIT_17 of inst : label is "B47EC40443F7F7047D0905AB665FAF513131A0456346BB6E9BD7A03D40A1C1E0";
    attribute INIT_18 of inst : label is "79A2A0D518DC418628E1C04CB2C307D859A2CA3D819B56AD5A51608B25805608";
    attribute INIT_19 of inst : label is "5FF7FFD1AF45555850A9F22361D7D785A803AB4447AEBFFC44410104115756CE";
    attribute INIT_1A of inst : label is "0E037E9A64C4CA8D47546D549173DCF7688BD896A5AFA3711BACFC44E473A96A";
    attribute INIT_1B of inst : label is "73BFB9A734E76D87DAB1FCEF3B1C270E378A0B1208F5833AF75AB5EBB669882E";
    attribute INIT_1C of inst : label is "C20A6D665454080AD886ADF2C801AD66B8D5C8F6FDAACFDDEBBBBDEF3F7DD7DA";
    attribute INIT_1D of inst : label is "51151013F7C7757B2CB2CB2EABEAEABEAEABEA9BB0B5DB6DA0EB1DE809BA414D";
    attribute INIT_1E of inst : label is "C510F090988A369088880D1498000083CEF3B3DD549DBDED4565467553CA2A34";
    attribute INIT_1F of inst : label is "0051005DAC708ABD6CF0406EA36DFEDBEF84C451B4577DEF7BDCDD5F73F28908";
    attribute INIT_20 of inst : label is "4A66A8F59AC93FC03050AB9D2DCF45BC05054447A8DB7412F856FB7B7B4DDC00";
    attribute INIT_21 of inst : label is "1062901090108D1AAADE3BC7A339EAEA0DE488888484ADD9D1D98484A1212848";
    attribute INIT_22 of inst : label is "2DB6DA51003BFEF1DE3B5476A8C8D0252202549A29C50002DE3BC76A8ED51990";
    attribute INIT_23 of inst : label is "4B51B788480C484C0868FACB6B7AF7AD9F7FFFFDB2CB2CB2E9252B30150174B0";
    attribute INIT_24 of inst : label is "2D71493264C99BDFA8801D9BD5CA7245F53D05ABD3CDEBB8153FE61991786128";
    attribute INIT_25 of inst : label is "C3E4755A05D8C3A1B600784BBB08FFF3E3F3F3F33A240005EEFE4666D9D4CE19";
    attribute INIT_26 of inst : label is "33B9D1B8CB107E77BBD8F2A2673B153843853843853868B22FF8BFE2F71D55E0";
    attribute INIT_27 of inst : label is "68EB5ADD6766D6A1BD1F93CDE4F37922A8EA730681F41EA024092806824ECC8B";
    attribute INIT_28 of inst : label is "A5652B329481A224458563B06760D23160306306738317FC18BDB53925C26731";
    attribute INIT_29 of inst : label is "29000002AAA80002AAA7935BB01B2185B3187CC0855CC3E7FBCFE1886BEC3DE9";
    attribute INIT_2A of inst : label is "4052024D2378B18CA9938BB815A41494DA0814C3A69B4D8C13AEBB18DA618D34";
    attribute INIT_2B of inst : label is "E9F6C5127CDCC5A1008A342001458045810AFDFEC89D37BF5580200D9BED8821";
    attribute INIT_2C of inst : label is "DE3DB501B52336532861B5320601DD8EDA626D6D20EF373068402281F6C512EE";
    attribute INIT_2D of inst : label is "C47189B9D69C15338B9CE2B7F1AE78BC3D453B52010C64D503571B41424C906C";
    attribute INIT_2E of inst : label is "24C9EE95B00552C4FF9627FC9C96C2CB2E660A05489DD65FEBA2A0F6B67E3D39";
    attribute INIT_2F of inst : label is "6EEEEEEEEBC3DEA0863287AAE2B9FDFFB0DE5E97D86F4BEC377CA5D4C8AAAD55";
    attribute INIT_30 of inst : label is "FFFEFA613DB002193A723864E9C8F3131296776443D9CE91BBD9DFC79E5DCB58";
    attribute INIT_31 of inst : label is "66CDF4554674546F40FA71A21439EF047A85EE05F93B32ADA6B43A567E79F7DF";
    attribute INIT_32 of inst : label is "016516EAAD8761A0ACF99FAA8ACEA8DD454D6C57057EFEADD77BCEACAB24B9B3";
    attribute INIT_33 of inst : label is "2502809511DF6ABD3B546DFAB64A3A3B9FD7B5DAA3956BDCD9EFFFDB2CB2F700";
    attribute INIT_34 of inst : label is "5A8C8107E485DCCAEE75974400805EC0096A5B922D8E90B889AEE731CA75668D";
    attribute INIT_35 of inst : label is "AD04AD1689EAE1E5689AAF4D81C61C461C601C7192CBB1861DFFF9B268201A2F";
    attribute INIT_36 of inst : label is "D86D97CDE8AF6F4A7AF4A759D64039B4C638D8BDC4B38D27524EE49DC93B9104";
    attribute INIT_37 of inst : label is "6E4A245429554B6E4AB4440855426E738996D3091B57BB233334EF55B39BF056";
    attribute INIT_38 of inst : label is "3D6110FC965D72AF39730C262D3247298B5542554B6CAE332952AAD6C4085542";
    attribute INIT_39 of inst : label is "29FFBC30322166CEE7FBE9917E47D121004AA22504882641B4745F540C47970C";
    attribute INIT_3A of inst : label is "E96472BF65FEA9588A8DBDAB64A2C678E8CA7A8FF5675002B0447EEAEE74A3A3";
    attribute INIT_3B of inst : label is "6AE67634BBAA24E8CE7CF322F1D1D9D8FE645E747D46D2739C63BB57DFA4C0BC";
    attribute INIT_3C of inst : label is "746C3FCFA6407A01AEAAD55567F5636B332ABA092ED4BC9F69AB64A03DA66241";
    attribute INIT_3D of inst : label is "F7CAB7DF4E951B6DD56C94747E3DB1FAF6DEA8EDF615F6D928787DF615F6D928";
    attribute INIT_3E of inst : label is "46A902115902002223515ABFECFCFFD9F90241C13F000070D4372483A64AC466";
    attribute INIT_3F of inst : label is "105BDBFE7F6B3BE985656BBA7274B76A91C93E458E72E63DEF3CAC46C6A132AC";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "D7834A65834A6406070380C054ADD4A5B69A3B7E449124CC4000003899C92914";
    attribute INIT_01 of inst : label is "CE4604020100481294E912727292529D724A10A94914201307F3EEE74DCE804C";
    attribute INIT_02 of inst : label is "FCF94432000117200640002380C99A4CAC5E368476865A3422A28A0F34CB9428";
    attribute INIT_03 of inst : label is "48B6C964EA86A5AF7B0208249D9A0FFFD8C3103AFA4437FDFD5548D88B9C9309";
    attribute INIT_04 of inst : label is "201381DC0203040414801710236D033005608C0F349B641858272F81520A0196";
    attribute INIT_05 of inst : label is "9918430E8643A18B7A60BA48FAE29F0228028DF0B34F80005C89441AD38F00C7";
    attribute INIT_06 of inst : label is "27EC90DA0735220D1B24C8250040002505414118158641E01339C9ECB1A81001";
    attribute INIT_07 of inst : label is "3309FCF958728D0494681CC80B311571102B8E9D41B87E8D481D280DA59078B7";
    attribute INIT_08 of inst : label is "05103732F684250AB39E464D13F65B4B03265312A4006750601D050DAC08D2E7";
    attribute INIT_09 of inst : label is "D30874B57D5F487F231C8B006E50B6415310C216C8049338B7D95050A3426E99";
    attribute INIT_0A of inst : label is "50C4363949E1E9B83851F95A6979584618410618400731CA2E2109097B1A4094";
    attribute INIT_0B of inst : label is "8463A2249BB0B22707081DE061039C04A27781944E701081DE8C000B24141482";
    attribute INIT_0C of inst : label is "2E21B781E17015C4340A621A105054D6D148AEA1A408189312A0D41698DD418E";
    attribute INIT_0D of inst : label is "4E09C13827044A060E042AF840CCCB97C949E0001400F8A09AD4014FEA6F31CA";
    attribute INIT_0E of inst : label is "08825B9A0D2ED60606190DA40D986B2586A06A98A112CFF658DB632E5F0CAA3F";
    attribute INIT_0F of inst : label is "1740480A0002920B55043502D56C1106B7AC15200200042023DFDC138B409AD2";
    attribute INIT_10 of inst : label is "ED0805200520A76944330829DA412094DC01492004C8320C1959049051049B6E";
    attribute INIT_11 of inst : label is "02589CAF400EEDB184BD30F9C35C8C25C8C2031FF225CC1AE444464461060D0D";
    attribute INIT_12 of inst : label is "68C068C31636831616027005C7391A2E3280020EB5684E98141452602AAA8285";
    attribute INIT_13 of inst : label is "021CDC4011CC60AF6B45735823D8D58CD60116247209045B8129C06C6200B124";
    attribute INIT_14 of inst : label is "2CD087A1B5006D594F393CA4F381008062291014F8439BCA00C72710018E4F20";
    attribute INIT_15 of inst : label is "288590B0111487C8B4C9085A4010084448C516D38A2871471F8141B202544591";
    attribute INIT_16 of inst : label is "E55D150C91C168D808207D2D2B2B8F8CC6D002DD047D3CBF4FF7F3E4808B2144";
    attribute INIT_17 of inst : label is "0152500502826117602597D7F383ED8A32335288355D0D7520B6CCF62B45C9D2";
    attribute INIT_18 of inst : label is "FB14594E091CA0CA7000C4D5040002B8DD9A8E5E4200000000864D38493484B9";
    attribute INIT_19 of inst : label is "47FFFD3E161800022361D7D785E803AB4447AFFFFC444101041155151400B95F";
    attribute INIT_1A of inst : label is "BB10514DB8C8D1125C19B44EA64A508FA5F6E352842337BDBDCCD3AF71BB2528";
    attribute INIT_1B of inst : label is "A0735F3CC95CD69D339BA2388E877845689B7A6C927D832F45366D24AD9032CB";
    attribute INIT_1C of inst : label is "0B6413516A2A028A8443C94090004BAD2D785B6CBB3D833700E6E338CACF9E64";
    attribute INIT_1D of inst : label is "C406444478584480020020014C1304C5314C130004C8041052004784B0432D82";
    attribute INIT_1E of inst : label is "0E597931392CDA400808842A4800000B7B5AD7242A44CB2998A9BA90AD84C440";
    attribute INIT_1F of inst : label is "005D9BA4B15ED14C096494B8CDA4424023C9C966D2290421084040A10010D0EF";
    attribute INIT_20 of inst : label is "5C88007807328016ACB2DFA4D452A94C2928286A336900FFE129090909004000";
    attribute INIT_21 of inst : label is "769D7676767664201145C8995C4281159451111115D5C44A4A4215D5C575715D";
    attribute INIT_22 of inst : label is "F4D34C0D3481222644C98A93111B2CDAECCDABC902A0579744C89931126AA376";
    attribute INIT_23 of inst : label is "8066D34202420246062356ADDAF7BD6ABCB37EE60020020000007006DA6DD806";
    attribute INIT_24 of inst : label is "7408100000000000E2800C201B749CDB7A441100A48780AD3A405C771ADD4E0C";
    attribute INIT_25 of inst : label is "BC1F670D394A8E0898D3B2B0506E3E0A180A180A1548B2CCD415204171F20F40";
    attribute INIT_26 of inst : label is "3BE832E23CA6BEE4F44AE1B40C2366817837816836818F06D95B656D855CDC34";
    attribute INIT_27 of inst : label is "88863144152B430897930D96C164B0CD8621E0683219BA6A4652337653201093";
    attribute INIT_28 of inst : label is "0E00700A4A92CCC08DB4B8B6156D1BB6650C36594C420F62107D82524A064229";
    attribute INIT_29 of inst : label is "E73000000002AAAAAA80A9EBC32B461E562100998CC86E4408881691840D0602";
    attribute INIT_2A of inst : label is "480602EB9828006C1B3403C0B1E22490A89D78CE106C20252E18405B8C09B8BD";
    attribute INIT_2B of inst : label is "5812CC6618818E0869F8C10D2F0934FCA44A01D490AA54800C2000020D841117";
    attribute INIT_2C of inst : label is "0A0018CA0847C281134C18D134F294A8202588A846962022821A5E1812CC2609";
    attribute INIT_2D of inst : label is "0A5211228B21860BC442E649A4F2C380C40C650CD35CC80014003E17D910A542";
    attribute INIT_2E of inst : label is "423159F65B34A0582402C1222A219190D198B46D228E619FE6CDCDDB81B56A20";
    attribute INIT_2F of inst : label is "A0A0A0A08893A219AE66A4BC2F0BEFC42941C03234A019085001503892900200";
    attribute INIT_30 of inst : label is "41020844FF2EEE14204428508110822220041200A4010002022B28F640E29104";
    attribute INIT_31 of inst : label is "10201989B8B988815416B7F964CBE0B49398ABB88B00CA60040129D4C1040820";
    attribute INIT_32 of inst : label is "B28C311865BD6E36B6D40933337311018A2B98DF34FC99C96192B51532DB6408";
    attribute INIT_33 of inst : label is "B73B365A3A00845E4D19B4484C3254CD2938C64C444E4B57F495EE600200104A";
    attribute INIT_34 of inst : label is "9731188A8A0A32B4194825BA6508A0400EBF65ADC8724F2703FCA4846FCE2A75";
    attribute INIT_35 of inst : label is "12891289120D9658912006105CE2CA63CA2CCA3CE1964CA3CE20C2050950A851";
    attribute INIT_36 of inst : label is "6A8B203657728091141B1004493EDE405747756E6A64B615282A5054A0A94289";
    attribute INIT_37 of inst : label is "80804BA912AE24808049A912AE24814A05494A922020D4C251C9D178C1501AB1";
    attribute INIT_38 of inst : label is "54CA72514C960CF472EA2A1554AA8B42D0AE04AE048242DD13255C090912AE24";
    attribute INIT_39 of inst : label is "D2816EA6A0B25D332A04171ADE151A1CA7B14B41950CA80A0280A02A201A7E95";
    attribute INIT_3A of inst : label is "8CCF4405892211A9D3368084C324B4935336A772CE43894543CE8A5C8DC3254C";
    attribute INIT_3B of inst : label is "5C2D93800CC4475316A52E35B51AA66945C6B6C6919B4A94A52ABD096CFB8D6F";
    attribute INIT_3C of inst : label is "A98953F79D0EA8E84B8D98E2C9664D804C0F43437C9AC1A82484C3240B4ABD00";
    attribute INIT_3D of inst : label is "0035402690666D10389864AB8952B592630311042CE2D330CC92A42CE2D330CC";
    attribute INIT_3E of inst : label is "8C906533A0E726744555F25FD7FD3FAFFA080404042449A23FC2CA5A918D4E80";
    attribute INIT_3F of inst : label is "A55DECAAB50056C16E198DCD5E38C7C9236F7ECC3994B64CEF69E18E8AA854F8";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "B4AA43A4AB43A19CCA65329966C966F84B65805C340D00623C00003859C8101C";
    attribute INIT_01 of inst : label is "034ED86D369B4DE0D4C90070708C189951839028460492803532826514CA204A";
    attribute INIT_02 of inst : label is "FC78143000050702860000A040C18A4C00423E6DA4C210F34C2010E6038DA1D2";
    attribute INIT_03 of inst : label is "00A092004283298B534A48C084502C209082103FAA44282AA2A02998CA9ABC01";
    attribute INIT_04 of inst : label is "100188C484001595942E185B3A090B4DA1142C0A241262A810020EB5522A9120";
    attribute INIT_05 of inst : label is "81FE2742A15028084CF2CC8773F16E508D5EA1F73846B8E30C3396D28293056B";
    attribute INIT_06 of inst : label is "49EC20060F3DCB6127024000000000801005028195DF0DE16AA947AEB022F336";
    attribute INIT_07 of inst : label is "BA81FC781470A9C0854C50C16599FB999CBD0F05002B5CF832D50AF661745225";
    attribute INIT_08 of inst : label is "FE5BB5E8F4866952A3AE868924F600420443598B9325E1CDE487154B0606D2A6";
    attribute INIT_09 of inst : label is "2DB15627566661450539A5CF921A497FD05BF7B248D34668B3D165F76CD90FFE";
    attribute INIT_0A of inst : label is "1AEC369918B1AD2C2978536708D3615869A61A618FE99E6F6BD23CCC96ECB2E9";
    attribute INIT_0B of inst : label is "8C49E77167307620802CB5108596A20030D040061A0820C351050D685756561A";
    attribute INIT_0C of inst : label is "6BD23F67674452679E2933CF3D5D56E7FCCBBF7977285A8B9AA2F597988FD127";
    attribute INIT_0D of inst : label is "5F9BF37E6FCE48B8B0B0F273E0EE6F9F4B86BA44844C5DB6F695A546FBC99E6F";
    attribute INIT_0E of inst : label is "2B8F129F1DA0B640C7D0E9BCAED6AB7EC0964AE6A15EDDF3ECC301BE7D08ABD5";
    attribute INIT_0F of inst : label is "A024048405149FF9D45155FE757C571E251CD4124125A5091E85581389E6F697";
    attribute INIT_10 of inst : label is "AF0474087002132450992284891858406C7448961A04010A283CB3CD2C96504E";
    attribute INIT_11 of inst : label is "4E1384AF42D4ECF69A1428784D5430D5434D3095F0C1426AA1A21A21A69A6A01";
    attribute INIT_12 of inst : label is "70F762EC14146C14144088139F7AC0DF1A132C9EB3CF6850954049429555A800";
    attribute INIT_13 of inst : label is "0D0C1CA04765CA1A2610D13086C993244CC2CC84602D01CD8E081FB62D3735D8";
    attribute INIT_14 of inst : label is "E8161B868705A1CFE3038C0E1128144A070380D099A183D6034317A806060E50";
    attribute INIT_15 of inst : label is "1DE33C62B8F09F5C70E89E386C542D00C5038CC30719F2060D1D4EB50628E3B8";
    attribute INIT_16 of inst : label is "A1515D4BC3C436503CE335CBE363E68FD98001B890008280F07807E901C778EF";
    attribute INIT_17 of inst : label is "0552000000EE76057382031E73632F66A0A118815D64CB2CCC97B13D9CC14550";
    attribute INIT_18 of inst : label is "5B04113710D44C09B8EC1250C323B0A8958A8E035816EDDBB690E18268842288";
    attribute INIT_19 of inst : label is "47D3E9045CB40007D785E803AB4447AFBFFC4501010411551514005451106857";
    attribute INIT_1A of inst : label is "37190BA6FE9EB99BBACCDBAEBD635ACBA28986D8C6B337B9BDC89840C3622508";
    attribute INIT_1B of inst : label is "CB6FC6BFFF9BF37A1C2F41D034B460746039D6769DA07EE520F1EB1B38F91AFF";
    attribute INIT_1C of inst : label is "1B2F1ACD2E2E2D555E2150111800B6ADBDAA5E7EEDC2683A3F4341D077835FFF";
    attribute INIT_1D of inst : label is "D73576F6DF0C7449A49269A5EEFBBEEBBAEEBB8916FCDBFDB2E94F8D9C612CE3";
    attribute INIT_1E of inst : label is "9F5ADDBDBDAEFFD88000077FE0000001AD6B57F73FE767ECCCEDDDDCFEFE6674";
    attribute INIT_1F of inst : label is "0045A8F10D3ED9F9A1E2D2FEEFFF77F9FEEDAD77FEBDCF7BDEF47CF3D1AE7F47";
    attribute INIT_20 of inst : label is "585504CC853A85D4DC325FB7FF3ADD78ACADADEFBBFFC477E33DDFDFDFC4FC00";
    attribute INIT_21 of inst : label is "45514545454543711132666D6626415133251515159587373737159585656159";
    attribute INIT_22 of inst : label is "7B64B7D554BAC99B3266CECD998AA8AAAA8AAA865E4BD08D32666CD999B33145";
    attribute INIT_23 of inst : label is "2F77FDD65216161212399CEEF79CF9CEBFD1A9879A49269A4C01548412414F94";
    attribute INIT_24 of inst : label is "702F75EFD6BD33335FDDDB7E1FF6D68DFB67BF9B37E39B7D3B66334CCF71ABED";
    attribute INIT_25 of inst : label is "5D7F74351B9AC66F2E11AA395B6AAAA8A8AAAAA89D402404C0610116E4F2A5D4";
    attribute INIT_26 of inst : label is "2A98B69E5EA0AAA7079AE3A40A1A44A84A84AA5AA5A8EB169EAA7AA9E15DD0F4";
    attribute INIT_27 of inst : label is "9C9CE7507E6D056F2A8A8556AB50A8C11E86EB09A0DC364F525AB864934C50C2";
    attribute INIT_28 of inst : label is "2A9150020080689C01243A24904803244161A8B08B44143A20A74A31E5269750";
    attribute INIT_29 of inst : label is "42100000000000000000A8821702121A56690053C9EA6263F0C7F338E6151B1B";
    attribute INIT_2A of inst : label is "40510067303009AD6172432411FC49848B870B8069A2C3000A69A1D03C390328";
    attribute INIT_2B of inst : label is "B4A080548555536F08528DE11A538469A012282AD11B711FB000000076580094";
    attribute INIT_2C of inst : label is "0C006B426B62D2D77B687BF3B610B9ADC784838346315515DBC23488A080148D";
    attribute INIT_2D of inst : label is "CC730CB2CFAE0790B4CAA3FF925282C6B045303E1159E23B84ED1770F35CBC80";
    attribute INIT_2E of inst : label is "42B8DBB7F8242B42475A123AA2A17170B55A860D0A9B3F9FE4A1A1FD95DD3A99";
    attribute INIT_2F of inst : label is "4A8A0B8B0FC9B078ACF262BFAFEFFBF5D896149ECC4A4F643C1F50BC5A85DBBB";
    attribute INIT_30 of inst : label is "B6CDB7873F6CEECD9B239B366C8E433330B2716CE6D9C5B3604B889014BCC11C";
    attribute INIT_31 of inst : label is "2E5C9DCDDDCCCCE4141C6D61445B24A41F1CCF3CDB114E3B636D1FDD26DB36D9";
    attribute INIT_32 of inst : label is "E26BAC575D004830A45D48BBBBB999C9DF6FDDCF046ACDEFBCDB9F9DBFECB397";
    attribute INIT_33 of inst : label is "8191939B3B37C532F45DFF6E675A9766E5BCE7766659B42A822A9979A49243C2";
    attribute INIT_34 of inst : label is "FD99D9DF1ECB3FD79FEF3EBE458CBFAFFAAA2F4EFC5E73F5C95EC694F1EBFE78";
    attribute INIT_35 of inst : label is "9B0D9B0D9B0FF7FCD9BABDBCCC20C330C30883082BFFEC20C35DA7974960B059";
    attribute INIT_36 of inst : label is "4BDE20FF7B9BEAD95EBF944D5B7AF6FE8563DDFB6EFFDC733AE635CCEB99D30D";
    attribute INIT_37 of inst : label is "E4EC6D8D1AE7C6E4EC6D8D1AE7C6E5AD9ECDFD9B793CF667E1F9972FE2106EC1";
    attribute INIT_38 of inst : label is "D9EF62E3DFFBCEDB4B9DB67B1FD8DE7B9EE7C6E7C6E47F741B35CF8D8D1AE7C6";
    attribute INIT_39 of inst : label is "2648B8DCDEB47DD99922FCCF749B8FE8E3F3E9FDA5CD2CCB32CCB32ECD9BA989";
    attribute INIT_3A of inst : label is "C4F5F89E348B99B9DBBFECE675A8D609D98B93B96F76F965728AC4DEC965A966";
    attribute INIT_3B of inst : label is "752ECDADD66675DDAB95999EFF8FB3332333DFE3C5DFF2D4A52851CCBF9E67BD";
    attribute INIT_3C of inst : label is "2EDFCBD7882BE0B8CDF7FFB3FCBF76C9E70594C9DEDCF13B0DE675A945DAF600";
    attribute INIT_3D of inst : label is "CCEECDFDBF777FCC9CCEB52CDFC920B8D3C999E717B3659D6D3F9717B3659D6D";
    attribute INIT_3E of inst : label is "F6854567B5456C76EC1DCA1A9DA9B53B53AFD7D7C46449BBFFC7DEE9BDEDCECC";
    attribute INIT_3F of inst : label is "F54B46AA25C14BD0BD39C6F975BDE5284C8D7CB34F57D46B9F911A35D839F6E4";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "6EBF4B26BF4B23DB67FEF239AABE0A8865D4C4AD3ACE9A3BADFFAA96CEEE7C9C";
    attribute INIT_01 of inst : label is "5DB8996A1BA9C98814140AEC2569E356A514DC04B4C08F775509140314274EF8";
    attribute INIT_02 of inst : label is "D3EE892D555D82998B9556933BBE65EB80572AAAFFCFAEAAFFE7AEAAFFCFA8AA";
    attribute INIT_03 of inst : label is "B445E79E34CC00242479B6906CEE6E8AC5D7BA80FF118228F5FDA45D32DEE7DC";
    attribute INIT_04 of inst : label is "7071A88A8E07B9B901E74CD9E6FA1C599ABE7D90EBB9D8EDBEB2849A9FBF9269";
    attribute INIT_05 of inst : label is "4DE7C481F31D4F17BC75829A37F7A08A57EE7CB62CB52CB21358AE80035AAA88";
    attribute INIT_06 of inst : label is "FB5B49A1D3EA497AFFFFAAAAFFFFAAAAFFFFD5DC07BF44350BB2233A13F67922";
    attribute INIT_07 of inst : label is "B4E12A56DF45FE446DD31C30ADEEBBBB8C927287314713B03E720E119DA10560";
    attribute INIT_08 of inst : label is "30C108DE39BC504A94E39BA6EF5BA6A6FABFAAF9D74C9AA46D6AAAA5599EB01C";
    attribute INIT_09 of inst : label is "65D744550324428A5DEF23FAD10ABAE0CC49D1F835DB720875806A21AD3A0228";
    attribute INIT_0A of inst : label is "A5AB02689AFD07267B06A2B1FEA4B31A10611A6145E2FEA2B5F8E4EEC6D7BA49";
    attribute INIT_0B of inst : label is "DD005A88A730A8A8420C8AEA290782AA30D4AA0A1DF4AA28510FA88AAFCEA74B";
    attribute INIT_0C of inst : label is "B5F82877FF94E7B869591A69D525AAB39D15199AF994E279C1E6B9A905FB96A8";
    attribute INIT_0D of inst : label is "D59E3EC07ACEE678F0F38000FBBBE3BF4A8CE528C07B3A0CF8772AC283D0FCEA";
    attribute INIT_0E of inst : label is "59A71E86FC506E6959F7E04D1956039E4FE5E87674DDE7F9D47DA99E97D7A195";
    attribute INIT_0F of inst : label is "5655A820679C4DFC767990FFDDFCA6593D14A9A061F70FDAEEB1300FCF517E00";
    attribute INIT_10 of inst : label is "47A6971D6C2615E5A9AA3745AE8AD056A5785C49DE82D47422E36104EBA61D73";
    attribute INIT_11 of inst : label is "50FCB375711BA387D1FEF6DEF396A8B464B305FF1938BF770D389FB914536E8C";
    attribute INIT_12 of inst : label is "AAAAF5554B4AD51C4A94F405AAAE555FAAEA4557A2BAC5D1D55575C5AAAA0000";
    attribute INIT_13 of inst : label is "D29781BFA6A93BE7B2A938CEB2AC64FC8BAAF3CF4802867A72F9D2CA53CAB5FE";
    attribute INIT_14 of inst : label is "28F6E5B93EF95452EF8F53D1F8EB7BD5C28E560A81BD5DBAFCC58AD1867456E6";
    attribute INIT_15 of inst : label is "BEA8FD23E2640839F89258FE9A7A7CD8E2AEBF95E2BA219EB2EA5EF6A2F2EFFB";
    attribute INIT_16 of inst : label is "0ED284F1A6925475C92408D53ABA3EA4087501DDAFD6694AA52DA5E5D6AECD55";
    attribute INIT_17 of inst : label is "AFA37FFF5AD247FF048EBD2662EA8F1688A8673089623BECBB90ACBCB3C7BDBF";
    attribute INIT_18 of inst : label is "2CBE49290B8E6D995FBB9693BA7E3668173DAD3FE3878A22466994CCEABEFD55";
    attribute INIT_19 of inst : label is "1436B0C5F2B2FFF756EFBBB8AFBB03BABEAAFAEEBBBAEBFFEAFEEEEFAAA89935";
    attribute INIT_1A of inst : label is "EBDD7ED50323A724AA2226D60D9394A362A9EEDEC9B12BB50FF3B6FE2348ADCA";
    attribute INIT_1B of inst : label is "1D67BADECB59EA2BB1C09DC79F3BD9C363FF39873082082C3A55007CA6B01F60";
    attribute INIT_1C of inst : label is "E38C62B08282275F2AAC9EA77D765B1C8FFA9E65039EA3B53858B66DB0442E45";
    attribute INIT_1D of inst : label is "A262AB2A23802C94AAEA2413CC33BF6F30CCFDF46FC1A288DA368C0B39CBABD2";
    attribute INIT_1E of inst : label is "80A1F810CB8E114FAA8AF6D29FEF32F1C1F0874683B84B092202B99B0E1E5554";
    attribute INIT_1F of inst : label is "5A2A27E8A082EEAE4B148B87CC308184B6813ACECB00389A8C2301EE8F6CC878";
    attribute INIT_20 of inst : label is "E011516517276CFADBE7B919A76566AD3D3DA5A766796E0E5E7DFA5AD9E49F5F";
    attribute INIT_21 of inst : label is "1111EAAA5111E88B51DBE622BB6DABFF7DB7AAAA04846888D5D5AA6A91219AA6";
    attribute INIT_22 of inst : label is "A34DB260A1584E917098E465662C2A02B1302ABB0459E86A7098465E263F1148";
    attribute INIT_23 of inst : label is "495DA3A89797282897ECF80F25093780FD448A68977982006560FF89155123AB";
    attribute INIT_24 of inst : label is "A1597B76CD53999942AAAD187E697B665F9F11E9F8C76918FF957E3F7F97F9BA";
    attribute INIT_25 of inst : label is "953FE18ED2940122E70DEA78C9D994E77676E7E5E47371C39C55AA8AFA30952F";
    attribute INIT_26 of inst : label is "1B958718E5EF4006ABA5E669DFC9985EFD6F5E856FD67AB9AE8EBA9AFFD5647A";
    attribute INIT_27 of inst : label is "DF6812865A506B22E2D4F283399DFD3EEE3BB000EC6708F1DC06AF231896A566";
    attribute INIT_28 of inst : label is "3DDA37932CCB79A6FF6346998FDB6198DBDF28A2DFC70ABA38FFAA2AFFF6AB28";
    attribute INIT_29 of inst : label is "10C5ABFE1111ABFE1133B87A51C380BE96401CBA9D45993964F8DBBEF78213C9";
    attribute INIT_2A of inst : label is "B83B80AAF07BA8A8FFF7A2AA33FE2AC0F4EA816008205110F3088BAE915AE192";
    attribute INIT_2B of inst : label is "EAFCA11B27AF8022D40F223ED076F8025941F5D64A26800054408AAA9A68EEB0";
    attribute INIT_2C of inst : label is "1ED521A019BA081D7A5121B7A5AE8B0D201F515123B38B88C2FFA0EE5E7D8BA7";
    attribute INIT_2D of inst : label is "CE737E0875EE380563FF1883EC5937431A77B9890C37518040CC0E6040BF08AA";
    attribute INIT_2E of inst : label is "8447FE39D6DB11A671378E9D1C1C70794CF56B80E2AD26E01F1A7A2E4CE71A89";
    attribute INIT_2F of inst : label is "EFCF4666CFCC3D275BB39CECC0BF8BA8A18E4349D0CFE61866EF3D809B6A8800";
    attribute INIT_30 of inst : label is "823B2546691A4440F2028102C80B18A8E8821048A6180922E5BACE2F19FBC5C4";
    attribute INIT_31 of inst : label is "DB83A223AAAA3112FBB616E38612532C35A1129F12F6B4184851466E0082CF3A";
    attribute INIT_32 of inst : label is "0862789CE99251F83C7AD275BBBB5551209A9B7E8601994993B80173B8F922A5";
    attribute INIT_33 of inst : label is "1FF73606886C9447D3A8AC67CC72A76BA028688BCC6D4122DD55E624AAEA2053";
    attribute INIT_34 of inst : label is "3BB85552E180779682E405F2FFC545550410D7B9E28F376598B98DEFE7E999A1";
    attribute INIT_35 of inst : label is "3183EE1A316C286B3315B16B4F3C0DD7B2C80D312CB231C7B3DD764B8FC4E0AA";
    attribute INIT_36 of inst : label is "FA214780FBB88DA43E2A49B28F157B19E2E3082C808F8841660BC906982C26B0";
    attribute INIT_37 of inst : label is "6DB3BB9BF2430B92B3C69B2D433C92A6E22FCEFEAB30676C9652E77001A27DBE";
    attribute INIT_38 of inst : label is "D8E854D4CE399DE6EE2231D13BAE1964B6C9A1163E6562237F0B265000FA16A1";
    attribute INIT_39 of inst : label is "1A01CAEB8D1C71DA68012ADED428DE74600FB720970F8B0E200BECF8049472AA";
    attribute INIT_3A of inst : label is "FC73516C301B77CEFBB84FDCE78619E5BB8C4772E922A061E0820954BAE771DC";
    attribute INIT_3B of inst : label is "49C8AA33640CE49D148786EBA82008C38488BC771283C8AE322C16206C6ABAC7";
    attribute INIT_3C of inst : label is "223161D7E7B0FC5D8AEE9A66E181D4962A70F72DB9A3BB7FECEED271B3FE9956";
    attribute INIT_3D of inst : label is "888579E035EAEB0B2A8BA58290269B063B30FFC04C8A789EC714A88F8AC79E35";
    attribute INIT_3E of inst : label is "3538595508BEC0B0EF8AA39032032046F8A25848BE0F1027947EB224333F7719";
    attribute INIT_3F of inst : label is "0AB43201BC8E0C688E023766F0493A20683CEA19911C3B7190F8AD93A0CAE662";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "13C0A0D3C080C6170B95CAE165CBE7F412030046609837A41600003890851213";
    attribute INIT_01 of inst : label is "045692492492581A8368A40A0A33546D0A6A4DA119552A81AAC27584EB09CB80";
    attribute INIT_02 of inst : label is "0285150A000858A2A940014844285F02FFD840204C007404C4022409C4044849";
    attribute INIT_03 of inst : label is "085B6DB6B245292A51A9A880949084209082102AAA4420A8A8AA0990A2D84002";
    attribute INIT_04 of inst : label is "7062251088042525164916B0C5B592000D28170335C214048025AB49444A2122";
    attribute INIT_05 of inst : label is "8C30260402010099400180184C0C8912F1100524114124921E492C1ADE000480";
    attribute INIT_06 of inst : label is "6C1280DA167416150000000000000000000061053D11E90F5A24401428AE8254";
    attribute INIT_07 of inst : label is "01020285080A4DC4926C142A5219999DD8E1004A22B27C480418201988511906";
    attribute INIT_08 of inst : label is "04B0A604A49498F10134D4C936095B50000319801309220D2808515C16B0C8B6";
    attribute INIT_09 of inst : label is "DA2C20A5551B0A40B090D2086C51248106B0421B690D98A28A531A0102042A48";
    attribute INIT_0A of inst : label is "3B1C8E4D63F2109CC240801838001A50410492490097ABE6E5638683534004B4";
    attribute INIT_0B of inst : label is "1445A0AA1C00A07BDF658A7BECB14F7D9629EFB2C53DF658A4880104110091C4";
    attribute INIT_0C of inst : label is "E563BB85B0209861164C308BF258466B6E62B33536249480D09C42128EAC5D16";
    attribute INIT_0D of inst : label is "0710E21C438840484A4B050418EE6C582C300840000006A60492491ABA6FABE6";
    attribute INIT_0E of inst : label is "4A090340433BF081D231421601A0B8A0028ECA04240A2C0A00C7823160F32890";
    attribute INIT_0F of inst : label is "1D53AA708658C6A148659428520494900628092992984360280D583F85460490";
    attribute INIT_10 of inst : label is "AF1448184C10260981304C09C24368988D5C326502380E0248DB4D36DB4DADAF";
    attribute INIT_11 of inst : label is "CA7297A830B10135161C32058A12ACB02A8B21300AB12C5815495495651602B1";
    attribute INIT_12 of inst : label is "C990D9A20021A20021BF3DF620C343A0E8BCE0E144A08F1E555591690000FFFF";
    attribute INIT_13 of inst : label is "0B1C9EC004E1382709C1384E09826486121B53434A487611AB01DB6C4A0D0364";
    attribute INIT_14 of inst : label is "1C70D3349E69271387121C487030184C040A0017816393DB02C737B0050E4F60";
    attribute INIT_15 of inst : label is "2D25A4A3A1045450A044D05048214EF42E7613C1AC237243583AEC74B1618461";
    attribute INIT_16 of inst : label is "144D955980009A8428A0758DA9298C4DE2F00E614FFDFE3F8FA7FC0D810A4949";
    attribute INIT_17 of inst : label is "090D550558CB41F0C2249D120A43998A0A0B923F210C8DB4888CC666295C280A";
    attribute INIT_18 of inst : label is "CD555D5EE702A0EAF702E596089C822F8531A1406844A952A4830790131C0C10";
    attribute INIT_19 of inst : label is "841A0E2AE1DC000447AFFFFC450101051155141400545111104141405401AF50";
    attribute INIT_1A of inst : label is "05B211D26C8C19DBC2CEDB8836A42B0A57563BA91AC25C2AA12022FE15C4D614";
    attribute INIT_1B of inst : label is "484DC4A7649376921BD24310C453D853D891623C9DF7DF4548FFE15B399E726F";
    attribute INIT_1C of inst : label is "192518590D0DE7F559095A219F546EE9B5AF5336CDB6E01A1B434210C38253B2";
    attribute INIT_1D of inst : label is "773774D41EAD01F1451C71C46F9BE6F9BE6F9B9126E8CDA498A26184946124A3";
    attribute INIT_1E of inst : label is "8F11D1F1F9E76DE2202207AE47EFCD25AD6B74B72E4793C0CCECCCDCB8F67674";
    attribute INIT_1F of inst : label is "CCC91CB24124197949E4D0F876DC77F1668FCD3B6F2DCFFFFFFCF4B3F2C61B87";
    attribute INIT_20 of inst : label is "4D00410D15A8C804140F58375F1ACC796D2C2C0E1DB70006052C9FFFFFC8F4CC";
    attribute INIT_21 of inst : label is "10401010101003300439672C66084000E38E044444C4C733333304C4C131344C";
    attribute INIT_22 of inst : label is "7A4804883E2811C338670ECE1988802022020087D03A338239672CE5D9CBB110";
    attribute INIT_23 of inst : label is "823B6D018181818181BBBDE6739CC9CFA2D1020F1451C71C5022D10B6AB68026";
    attribute INIT_24 of inst : label is "C64A80000000333382A000B20D9B5E1D8DA7457F5A083F320DA882288B713360";
    attribute INIT_25 of inst : label is "957C17A10800005A00701094302C2A0818080A0AF1200092D02044C016C27498";
    attribute INIT_26 of inst : label is "A225202094A3AAA050200530446066D26D26D06D06D00D26C0AB02AC11429E2C";
    attribute INIT_27 of inst : label is "C614A5060001605A02910A8542A55227D03425393048E16F5E5A51C46828901A";
    attribute INIT_28 of inst : label is "4A2251084A1202015031AA06940D2E060C79E78EF0040980204C886A9290C961";
    attribute INIT_29 of inst : label is "C6300000000000000001B7801A800A8B55FDA80563BCC7015E02BC4210570853";
    attribute INIT_2A of inst : label is "1FFFBE8C6F09A45116852CD2A61C6E1580822A2A490492012A412251294D12A8";
    attribute INIT_2B of inst : label is "56542B0488A8825A38000B4700001C100401282AFF6361558A60001C00905506";
    attribute INIT_2C of inst : label is "C2564A404A4062E195064A4D50500001049032B24E022A60168E202E542B4490";
    attribute INIT_2D of inst : label is "18C4203AE818071DC3201505B6580020060245AC700A8B2A80AA018295522F93";
    attribute INIT_2E of inst : label is "C810050A018182CCF11667892920303040B1952877418A5FE04547FDD019B30A";
    attribute INIT_2F of inst : label is "25454464401D4358054460D13440202046094B402325A01381824920003552AA";
    attribute INIT_30 of inst : label is "3CD9E634C08555020C0C04083020166647388C79BCF331C4458A280808001CA7";
    attribute INIT_31 of inst : label is "30609DCCCCCCEEC59A1CFB1071FA14319D698D49BA9250FA404901AA0CF3679B";
    attribute INIT_32 of inst : label is "2ECA29B4D0140C223770823BB9999989CBA1CE80A1AA0C21891B279D9F734418";
    attribute INIT_33 of inst : label is "921D7AC32362EE85698EDBCE66584669071CE778666755FDFDF5E2F1451C5800";
    attribute INIT_34 of inst : label is "F99B19982F5B38C11C62663CED99BEBAAEBAAC5EFE655BF6360238424DE09F7A";
    attribute INIT_35 of inst : label is "9B6D9BED9B06D7FED9BEF158A51040940106004106FFE004117E3B1B3B69B4DB";
    attribute INIT_36 of inst : label is "CACE36747BBBC5F99E5F99FE7FBAC5FDE8E3FDC29E3F96FA6DF4DBA9B75267ED";
    attribute INIT_37 of inst : label is "C5996C8C1EE0A6C5996C8C1EE0A6C52160AD815B3108E66B26DDB3A28CAB21C1";
    attribute INIT_38 of inst : label is "C277EE05E7D88EBF6ED94582D816CE93A4E086E086C4165C183DC10DCC9EE086";
    attribute INIT_39 of inst : label is "9072301416A2819A41C8588B60928B7283C9606D11E88CFB3ECFB3ED36180D61";
    attribute INIT_3A of inst : label is "460865B14833983119DB6AE66585006199B613BC610C230C7658D18200758466";
    attribute INIT_3B of inst : label is "172BC3CDC8866399A615C116C28B33482822D822D8EDB8CA729EFDCE464C45B2";
    attribute INIT_3C of inst : label is "8CDB080849CA2EA150FFE2337E39171BC0901376021E512A96E6658611FACE00";
    attribute INIT_3D of inst : label is "CCEFD8B15A43B6E09CCCB08CD30CB5BF178A19D74633759968B61746B3759968";
    attribute INIT_3E of inst : label is "D83314AA3314B64675A010CA99A995335348646404FDE9822BC0EF61990188CC";
    attribute INIT_3F of inst : label is "B04C76FE51D263204658C6ED1CAD64436B728219A996C47D90684D1CEB473608";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "2137E5E43736E7979DA1F37955D4C00D8E30C521531490556B555585BC419C44";
    attribute INIT_01 of inst : label is "5463C40CE9662C1F8B3AF16F321804B8531E7BF41C9555444646F3D95919D3C4";
    attribute INIT_02 of inst : label is "D561CC1455518D59F055A9F1F1C05A353F5F5F45745FD47DCFF5D47775DDDD55";
    attribute INIT_03 of inst : label is "5D163CF3BF95FE7FD965F0CF1B915975C5D7457FFF11755577777C84BFDF25C1";
    attribute INIT_04 of inst : label is "5517FDDD54539696A5701449D9457D5D2DD31051175415E575CE56744737B36D";
    attribute INIT_05 of inst : label is "97141E7CC5C7146C555474575151D55545A71001E15FB6DB375C10FFB7F48145";
    attribute INIT_06 of inst : label is "C45D4535A975F9B151555555555555555575A9EEB54EADCAF4C47DE7174DCBFA";
    attribute INIT_07 of inst : label is "D0152B9C79D652BF147DE23D5A5544441165CC6B6596ED17ED98F56EBF4DA2CF";
    attribute INIT_08 of inst : label is "EF0CED3F967BF429499659671DD874764DC4EADD6CFBD1B6DB97BDEBDE355DB3";
    attribute INIT_09 of inst : label is "D3641EE3FD8EEB00710E0D652479C30467262F8E7F64EFDF7DD44F0EA362FD55";
    attribute INIT_0A of inst : label is "7D50D52355C55C1554794F33D1DF316CB6FB2CBADF398F3B76C6F9C7BBF3FFE9";
    attribute INIT_0B of inst : label is "F654E557055F55177FF71510FF7D5D00DF544004F5770041517D05555989E187";
    attribute INIT_0C of inst : label is "76C67C7759B35A3286B65CF56E9CE7257384DD5146675B461C254729E45DCC15";
    attribute INIT_0D of inst : label is "4664115E911714588D8F555549551D052471BBC515318133159E0E7FBC395419";
    attribute INIT_0E of inst : label is "A4D34DDF649453CA6ED93FFE4B597ECF1D04A0DB4679B0ACF1D7D9DB68104381";
    attribute INIT_0F of inst : label is "54D565554D36C75054D320545563E18667D754154D55526963DF8BCA9F5E40FB";
    attribute INIT_10 of inst : label is "7A8783DCFCA0751DBAA8D555BAAA1754ADFCB4493FA49E78EBAE4596AEBE997A";
    attribute INIT_11 of inst : label is "ADA3A917DADA51E9B8BCF2CAC708DB6E81C6F7BF00601E9A5BAFA68AAEBA9E21";
    attribute INIT_12 of inst : label is "BA8A4555AAAA55F5AA8A77FDAEBA7555A2AB55558AAA4775EAAA4555AAAAFFFF";
    attribute INIT_13 of inst : label is "A762BCDB6AA2FDFFEABAFDFF2ABAFBFF2AA8FFF495E6171E262EFF58A612FFBF";
    attribute INIT_14 of inst : label is "A9AFF7BDEACE65D3FA0B15D0A0BEF1D0A10B178D1F81F5B029D84BD59E06F6CF";
    attribute INIT_15 of inst : label is "185AA17C7EEDB69561A154BAAAD39DC2C1932EFF91193DEF428669BD83BA8BA2";
    attribute INIT_16 of inst : label is "F2D89CC06AAA45559C71139170781E7190CAF557AFEA7D4FA2AEF515EA46C951";
    attribute INIT_17 of inst : label is "9E83BFFFABE7D8263B18AD7AE7846DDF5554F7580AC3ADF766B3C8B706BA0823";
    attribute INIT_18 of inst : label is "88EB5D0BBAA8DB380AA42590CFAA6C7CB268B276C63ABB76BAB1C51D86E8D591";
    attribute INIT_19 of inst : label is "680008BFFE16FFFEFFBEEBFFFEFBEEEFEBEBBFABABFFFFFEFFFFABFFAAAA43A7";
    attribute INIT_1A of inst : label is "AE997D75C6E69506CE66165435E0AF6340021B2D1E05473FEEEE8555C9F95AF6";
    attribute INIT_1B of inst : label is "7BFA0B78A6FE859CECE6776DB1165F8A47BB30FD2A80FF7A255514E712E9B79C";
    attribute INIT_1C of inst : label is "EFBCD0310E0E45552AAEFE872AAB5BF99ECBD36566CA93176919E138B19416E5";
    attribute INIT_1D of inst : label is "80027557E7089DC39618E79DAAAA1986AAAA666798E45965F0E9A47DF8BF7DEF";
    attribute INIT_1E of inst : label is "8B869038EFAB1967AAAA76598C98455DA4A9F7E62E89997166469999BA6A455F";
    attribute INIT_1F of inst : label is "AABAA9F5B8E1E797EA8AEDC9BE697E73E9ACDEF7A7A6D7615A967DF5599BE7AE";
    attribute INIT_20 of inst : label is "594414F5FD7C2EA46F5E4BDD1CDB56E1B0F094D7D8C7675248F35B7B0F11D7AF";
    attribute INIT_21 of inst : label is "77EE5111B7775775EE6910FD54115511F69B4000D595177766664404B5650040";
    attribute INIT_22 of inst : label is "3E7192E4C14F5EBDCA6FF775DDF72982DDDD2A1A7D361D4CCA6FD75CDBE45551";
    attribute INIT_23 of inst : label is "A6641C15D5F51515D59503F05ED7D83EE3AA08CF24963CB385740CFF5E65C432";
    attribute INIT_24 of inst : label is "28B62B76388CDDDD375F08D291F76354A46C11CD4797CD51346AB75DDC6DE5A2";
    attribute INIT_25 of inst : label is "961C6E90774FFC09C857061766476B5C99995C5CF565CF3E95554555D3E7A81C";
    attribute INIT_26 of inst : label is "4C6ED43E373D400E5EA4B1FD6EC4DD3FD29D3FD39D297995FBF3309CBD6332CF";
    attribute INIT_27 of inst : label is "D53760321D3B2409C79246FC85E70470E779A9FC1611E6266E9994F9D479C443";
    attribute INIT_28 of inst : label is "B7460C59739CBBE7759B647D7D67567D6DDF55555D5515DE5575575955F77451";
    attribute INIT_29 of inst : label is "E775BBBB5401BBBB5405F1E33DB6F98AB5D6D7C1FF7DD31105985F83B41DF743";
    attribute INIT_2A of inst : label is "317100475755FD5DD5F54754573555556F15D0D0BEFF612DD5B6A97D6BB1D313";
    attribute INIT_2B of inst : label is "C495FEF15191FB09797C04507F1B43F9E5535201AB661F35553F10156927661F";
    attribute INIT_2C of inst : label is "D558B3F4F6E56BCA44B0B3EC4A7D294EDB5DE343705CFBFC3D3413D6BD17CF3C";
    attribute INIT_2D of inst : label is "719C14779971C3BADF46F134927FD4EBC31CB8915749BE1995BAE0CFD46635D6";
    attribute INIT_2E of inst : label is "E1294BECF1537AB50E9072BEDED76667B31BCDD4DFDBCE0AFEE7B1AD67185FB4";
    attribute INIT_2F of inst : label is "19792525789F7A1CF467719430CC3D332F30AEAC3339E4EED0B10D6796170199";
    attribute INIT_30 of inst : label is "9A6E44B540E257B331BE6ECDC6F884441A9F9C596E7F796490C9286E26349CB3";
    attribute INIT_31 of inst : label is "AC6E7FFF6666FFCC2868D6EB04118DA568B0FEBFD1199EA7BAAE536EBA6979E7";
    attribute INIT_32 of inst : label is "2BE1F191BAE8C786682A9255AAAA55314B2699D72CBE18318E693151A9AE646C";
    attribute INIT_33 of inst : label is "E1BB3E9FA9BEFFE4BC66E7D9BA2F99996EE69F79ABC2F7DF2A00F7778618C79F";
    attribute INIT_34 of inst : label is "6AEF7774CEAB1583C7A34559E6AB6FEAFEBFFE75A5EE1D6396FA31C4D2A09917";
    attribute INIT_35 of inst : label is "F92EF71EF9EAEF9DEF9FA928C4922449492424929A699659082A7739C1B4F067";
    attribute INIT_36 of inst : label is "A8E65624EAAC9997FBE679969AFFA559CAB257F30E9A02413A4ED907E93A66D1";
    attribute INIT_37 of inst : label is "566ADEDFBA6AEDCD6AE6DFB56AEECDD5AF8E15BF95AE999FB6F26CFFB002D5FC";
    attribute INIT_38 of inst : label is "ABA35C9DBAE89496B93B514169389A367A6891B5EED6340C39BE4331EF38B5B1";
    attribute INIT_39 of inst : label is "AEFF76DABA7196669BFFE37FAB0FFF97826B979DEE9CFDCF9A67F77C04735533";
    attribute INIT_3A of inst : label is "2C1B4D699CFE5764EAFB4954AADA1961AAFB4556A0E46651AE28994366AA0D54";
    attribute INIT_3B of inst : label is "E084D6DEBFEA9E66E9BE55B94D09FF59FFE2E17F666E7BCF2B4AFDFE9B246E73";
    attribute INIT_3C of inst : label is "E66743CF232A9E7F06AAB666AF988516FF003343FA6649A63BAB5D0C66AAC55E";
    attribute INIT_3D of inst : label is "666F9F792F3979F0E666F5FF67BBEBABE2CF660F9A999A66BC69D75999A2669D";
    attribute INIT_3E of inst : label is "5669515D39AE4104FB2A605AEBFE356DAB1AB4B43EF602EBAAB9FB44E66E7599";
    attribute INIT_3F of inst : label is "9AAF49AB9649A72981E6D982D706989A949C424C4E7AF199605020CD648189F7";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "C0A00000A000011088442A15000000044B648024000009223E0000F67082181A";
    attribute INIT_01 of inst : label is "0B1CDA6C361B45F45247FF61650E8848E1D108108721BF8890130026004C2004";
    attribute INIT_02 of inst : label is "80500124000402002480008085972A3900077FEFF1CFC6FF1FE7C6FF8FCF8DFE";
    attribute INIT_03 of inst : label is "00249249200811C0754042C080F824209082102AAA442AAAAAAA9EB0C6885C00";
    attribute INIT_04 of inst : label is "7001FDDF8000B9B9E02D544B8A4898D920046601004309840001423400224800";
    attribute INIT_05 of inst : label is "00620040201008103EFE3EE3B8F8F777E2582006180030C3DC2892C1D61801EF";
    attribute INIT_06 of inst : label is "01090001DC74C9683323B45AB1AAAC5A8A089FC8F45B44B433384CA208184922";
    attribute INIT_07 of inst : label is "1D8080500C2160048B001D816588888C889300840103137C12C21651E1940900";
    attribute INIT_08 of inst : label is "964B30F2E626E0C13B8E0E0C00848000101188EBB924C024C480564487E041A2";
    attribute INIT_09 of inst : label is "24B921015501138E4435658B0002C965804B00000001282082413364C993036D";
    attribute INIT_0A of inst : label is "0A05028100B0040C031807030007031A61869A6182CD8A62214320E078FFDB59";
    attribute INIT_0B of inst : label is "0101899B6FB0F701C00C3C380187870030F0E0061E1C00C3C3870F782252C388";
    attribute INIT_0C of inst : label is "21438844046EE335D7719AEB9959E63165C39111163AC219095040AA290C1006";
    attribute INIT_0D of inst : label is "93526A4C4988B4202023800016222C587086A064824C429978C12C83E9058A62";
    attribute INIT_0E of inst : label is "634D184510E1B00A3B89E04D92041A122051AEFE1B2E850122820DB161EB03D5";
    attribute INIT_0F of inst : label is "F07E0FC032C9DFE0032C9DF80094C69A30BCF03F03F00CE13E857055080178C1";
    attribute INIT_10 of inst : label is "961F746370639C671CE338EF1BDC78F1657021B61F8C6307612C92CB24B2D247";
    attribute INIT_11 of inst : label is "260180A1D27842C61A1428424C1930C1930D101504D19268C9A61A6986187792";
    attribute INIT_12 of inst : label is "1E3F1E3F1E1E3F1E1E001C07C71BDE3F8FB1EF8E37EF0C1800001FEE3FFF0000";
    attribute INIT_13 of inst : label is "2C280E60738CE39C671CE338E719C7B8DEE3DF8AB166DBECAE0244B68D3FFC7F";
    attribute INIT_14 of inst : label is "8407886200C4802C6001800600180C06030180F585A509CD4B0A039896140730";
    attribute INIT_15 of inst : label is "30C618C659CCCF6CC0896E6008836100510998060331C404080C261302986619";
    attribute INIT_16 of inst : label is "C0CACB37F3C71EF8B4D3D8024848414610600BFDFA83C3E0F0780FEF82CD31A6";
    attribute INIT_17 of inst : label is "141B0000016D3728B90008508C8456C17574F0550283065B006B601B002B93A5";
    attribute INIT_18 of inst : label is "CFA288C4319900C62180C10C82860B0E8601E48980B244891211608724800200";
    attribute INIT_19 of inst : label is "0C1A0E005284000101051155141400545111104141405401550001555556E841";
    attribute INIT_1A of inst : label is "2C3903A6E4C4D8CB3646596B3108421EC00250C2108616E0B74CE15420738421";
    attribute INIT_1B of inst : label is "F7D9E9F66DF67B76D86EDCD73580C700C71118120800803D25FFFC5B3A5B082E";
    attribute INIT_1C of inst : label is "EDB69F04ACAC1AAA800741501FF56EA1B5E840B6CD86DCDADB5B5DD733B4FB36";
    attribute INIT_1D of inst : label is "88AAAAA92D0A2021045141062288A2288A228881BA20B24930DB89F6DA7DB6D3";
    attribute INIT_1E of inst : label is "8B286CC484832CB0002209AD85454501AD6B5039AD89658444644466B2C6222A";
    attribute INIT_1F of inst : label is "FF1286BF39615D6CA1A2626632CB9C91CB66661965AE794A52941EBE51935905";
    attribute INIT_20 of inst : label is "B455052DAD19A4C0B01B5439598E466CECACECAD8CB2E4151DAE725252429F00";
    attribute INIT_21 of inst : label is "CC000CCC0CCC19154092324623A6D400A92E77777B7B599191917B7B5EDED3B7";
    attribute INIT_22 of inst : label is "5B6DB2C014364C999332C66588A6038019B800330861000093326658CCB1940C";
    attribute INIT_23 of inst : label is "491965C1C1C1C1C1C1C89CE2739CC9CE80C5AA531045141068111014914925BA";
    attribute INIT_24 of inst : label is "5D63CB76EDDB99996AAAA438C5B6F3C58B79449B36525B367B73365D8B797B34";
    attribute INIT_25 of inst : label is "C1E5251201B84023720018090BA9EB323232323290092492FEFF67F77C8A2402";
    attribute INIT_26 of inst : label is "3B398338C7206A3359D840A4A733144A44A44A44A44A28B2AEAABAAAE5085440";
    attribute INIT_27 of inst : label is "7C4C63BC46E5C4237A9CA05028140A0098A62B04A1EC0C8444229886090EEC23";
    attribute INIT_28 of inst : label is "A201101806012024018878303060563060C30C30C3C71F1E38F8FF7BE3F6F079";
    attribute INIT_29 of inst : label is "4210141414141414142280234203034A1031FCC1A0D82367F2CFF18C63E519C9";
    attribute INIT_2A of inst : label is "000380EF807A3DE1F8F7E0FE307E7C55120003D269A6C3C00061AB381E658138";
    attribute INIT_2B of inst : label is "3B20D01E24E4C3230006246000C580038014FDAAD433615FFC4030109258A810";
    attribute INIT_2C of inst : label is "1E8D2101212242391125213912001B8586A061E10609393048C0018B20D01E24";
    attribute INIT_2D of inst : label is "842119B0C48401188009C8B7DBD278A63C44AB1201145691024710C0418910E0";
    attribute INIT_2E of inst : label is "3659D0A1208018C077C603BC80824041264200000AA52E9FCF20206622D9B330";
    attribute INIT_2F of inst : label is "6222222233A90A208A288795E57A1A1938C447049C63824E274C3584C9088911";
    attribute INIT_30 of inst : label is "9264925002808A1C38763870E1D8F99990972126464C8C999528577187BAAF4C";
    attribute INIT_31 of inst : label is "A448C44444446647005CEF51005816885918CD18D81B2C0926243EB27249924C";
    attribute INIT_32 of inst : label is "01671ECE398060510E5024888888888C6BA46C4840546D45AEDB5C8C8B6C9952";
    attribute INIT_33 of inst : label is "801102ABABBED00A74C65972361C22326DC6319623C22A8AAA80A43514107100";
    attribute INIT_34 of inst : label is "58CD88898D8BDAD5ED6BB6AC4D89B010055450A62D5C50B581504610C06AC658";
    attribute INIT_35 of inst : label is "CBA5CBA5CBE2C16E5CB54218818619165964596596DB6186182843164B74BADC";
    attribute INIT_36 of inst : label is "08EE01D9C88E42DEF32DEEDBB6C00865C078A2A52CB65136166C2CD859B0B125";
    attribute INIT_37 of inst : label is "C6D82C650ADAC2C6D82C650ADAC2C67B1D85FB0B11AE223373788F2B3880E0C3";
    attribute INIT_38 of inst : label is "1F6BA331B6DAE3D9DB332C761FB0C65B96DAC2DAC2C659430A15B5C5850ADAC2";
    attribute INIT_39 of inst : label is "26DCBCB8B371608CBB73DD8B6A160B2082C1656689944E7B9AE7B9AE245B7B8C";
    attribute INIT_3A of inst : label is "048561B201CC88B158CB302361C2C20888CBB8896A2EB3046608E5D44C61C223";
    attribute INIT_3B of inst : label is "3420FC6497622188C9BC9B16C40B11937362D882E46590F7BDED0244B606C5B1";
    attribute INIT_3C of inst : label is "446DDE1C630009000C22CB116CB232DB7F954821504454083B2361C025C21621";
    attribute INIT_3D of inst : label is "66456FB29D119658C46C384464DB4B41218D888196B161D8744BB996B161D874";
    attribute INIT_3E of inst : label is "500B04A2BB04B45723029C355D55EABAAB964B4B3A346DB595390DBB2E458AE6";
    attribute INIT_3F of inst : label is "B3A4A7AA126B0B238364622086A666709385C0D522F2DE33E071A956C603734C";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "DE09BE5B08EF586E414F8D06EA2FFF1363C73BA080605DAEFDAAFF23C401FBF1";
    attribute INIT_01 of inst : label is "014FBDE8720F1BB586CCAE761A5E555DBBE24C613F85CF913D07754E641EF111";
    attribute INIT_02 of inst : label is "D42332F5AAAE634E886AFF6E9EC655DD3BA3AAFAAFAFFBFFAAABEBFFE2EBF7FA";
    attribute INIT_03 of inst : label is "30885555600AC619759146A5D17C31759082457FAA4477770000C1D1A4C86016";
    attribute INIT_04 of inst : label is "EAA2BFFAA6AA070F3CB6ACB0722B75269B6D396EEDEBDF3E9A79750BF88A6CB2";
    attribute INIT_05 of inst : label is "C05742113159791964551151558159D9034AA50F9C6220920E018E9617A9FB14";
    attribute INIT_06 of inst : label is "3A5C3EDCE49EB4DFAA2AFFFFAAAAFFFFAE8A615636AF2BA3DB9CDBEEA891B299";
    attribute INIT_07 of inst : label is "15C32D9DCF5B6543DB8B1F583D88DD998EB49CCB524D4F7853E6269542A05535";
    attribute INIT_08 of inst : label is "79E5E42F8D999E5FB1FFF2F1E2D8DBDBB21F3732D79F0FCA5E6EEEBAED96F7DD";
    attribute INIT_09 of inst : label is "65DF15D403735847BC73AA989A122CA3AF4F545C209B19A2DA11B869DFFB4AAA";
    attribute INIT_0A of inst : label is "B8AFA9FEBA1BC3F3A5F6FDD226E9D0F19249F3CF6DF623DB4B509819B5972936";
    attribute INIT_0B of inst : label is "0D059A8A71104DF70540C41741045DFA00455FF91020EB7C0405F1D147471AA8";
    attribute INIT_0C of inst : label is "4B506418969539CA3D8566B465F50DC4CF6F2EECBD133D353BFEFE5001863FF9";
    attribute INIT_0D of inst : label is "C790660941CCC9AD7D7E05044A23705825A46523C14A758C29E521C81FCC8971";
    attribute INIT_0E of inst : label is "85F7D3EADA4AFDB5ADA62DB20897768FC27AD0BAB2FCA6ACEC6DF26B8A18D2BF";
    attribute INIT_0F of inst : label is "0014355570146F0C130116C344D51EFB5BA411D54004483890A4253E0D216D94";
    attribute INIT_10 of inst : label is "B4F1028CD7DD114435DA01846C4D00445BD3EC2074738AA4CD1004121044A9AF";
    attribute INIT_11 of inst : label is "4A4A14C11CB1061E77062D4160F1618118606071061FC3E5337179277DF7EEF7";
    attribute INIT_12 of inst : label is "F63C11704949301449D56001C46D102010554409E41940211555040400000000";
    attribute INIT_13 of inst : label is "419A1730D6490060B37500C0532C00409999200E67DDC8A1E34848A2618F0000";
    attribute INIT_14 of inst : label is "524C9224932A350144F556914E412A955CFD538FB35EEF61D0264FD06DFABD80";
    attribute INIT_15 of inst : label is "C307C85251D7FE601FD4622DDD59A0055ED18802DCC1805CCB5112020F132208";
    attribute INIT_16 of inst : label is "B1798084D4D50051021855D497172AD5CFD50310052B35554A8252485538A490";
    attribute INIT_17 of inst : label is "69077FFF54002F3CC2E71091597B360466679015A57F1288991C2658F914C3C0";
    attribute INIT_18 of inst : label is "8D51597E826197CBE3699ED41C6D56BDF920B6D429083154A98F55D15A13945D";
    attribute INIT_19 of inst : label is "143E1640B8ED000F56FE0101FAAA551454545451004041410104015514141009";
    attribute INIT_1A of inst : label is "02E05764A88A11169888964E6BBAD6AA78A28796B93A55BB7DDBB45186C0BD6B";
    attribute INIT_1B of inst : label is "B901FCB718007833B28B9CD7DBA9C3517B004B02D0222A98125AE918AE220863";
    attribute INIT_1C of inst : label is "5200D0F1484A07FF86419CB5655449016C3B87258B25939716B2F47DDACB1AA4";
    attribute INIT_1D of inst : label is "826089088A69A4243AE304025C57A669715C99A00399869AC43049A6898AA6D0";
    attribute INIT_1E of inst : label is "3240113160344964BB1946283D7722697A5EC0A65B12595988A988986DA0545E";
    attribute INIT_1F of inst : label is "FFB4B6883615597374159AB241908984B1986B0A1B78381A8C210A8E851D5895";
    attribute INIT_20 of inst : label is "FEBBBAA303736A3F9CBDA942F725BAC246461373271909FA5B04AC8CD9EE2955";
    attribute INIT_21 of inst : label is "5515A2225555B80B11D66692332DAEAECD6488C81555B884D1D1808045552808";
    attribute INIT_22 of inst : label is "F38F69161EF8A3067D981B8A222255D50888556CF3C7D73F7C9918A72613EBAA";
    attribute INIT_23 of inst : label is "C91B7281545085855048DD37318C0DD282C5FE22965910416881444523827285";
    attribute INIT_24 of inst : label is "A29134C946716666E00042CD6E780C3B23DFEE76BD7AB6E8A3D9896221828CC9";
    attribute INIT_25 of inst : label is "5148122181D915B8371868680FB594B96C7CA9B9A1121045C455985D4C4AA415";
    attribute INIT_26 of inst : label is "B952520A78E23F68A9F2E3B69D1F43236376233276378F06E60FCD6F73AA42BD";
    attribute INIT_27 of inst : label is "415DBBE0476100B830CC9594303839458922794AD866385BDC5439D248B7153E";
    attribute INIT_28 of inst : label is "082BEF66CCF38CC9C47123E4921C9DE41E28F7CF29EAFBBFAAAA2AEFF8AAEFFF";
    attribute INIT_29 of inst : label is "529A5555AAAA5555AAA3C6F4838546D6117185476FF405A3056C0883310154EF";
    attribute INIT_2A of inst : label is "12AEFFBEE6AA9FFDAA7BBB6BBBEAFEBFF86E6091924D286E4C9230D3F9813AC5";
    attribute INIT_2B of inst : label is "3A691A363F5FC8B88C436BE5997D95309444FEFF4F5134D4C000CFFFD7CCDD56";
    attribute INIT_2C of inst : label is "AAA282DED7F8CDC72FCA82F6FDB2E26369129A1AEDA52840F1C9FF34C3C44CC3";
    attribute INIT_2D of inst : label is "8C33EAC3594650486418B78AD39E63284D614424190D982AC1765DA495DB045E";
    attribute INIT_2E of inst : label is "C8366BE8FE2127D7AC63DFAA2B293E3E95783F744AB2EAEAE1DBCFC93FE26F4F";
    attribute INIT_2F of inst : label is "76363A3A227886B9965C22D6E4700C0A9DFEE262EE773E977F1863E9515DE8AA";
    attribute INIT_30 of inst : label is "61990502FC94824CE20599328807422261641048A59149227F9FAA962BF17112";
    attribute INIT_31 of inst : label is "5B818000B9BB2203559B5C55FEC5569C9A1F85018560727E878812802186C71A";
    attribute INIT_32 of inst : label is "BE1A38946207941A07F5791155511171964A89896EEA887949969515521800A5";
    attribute INIT_33 of inst : label is "8E4C02682E4D2FEC139998A6CDA6E66B0329608A5414FD7D5A0DD3043AE33600";
    attribute INIT_34 of inst : label is "B7133FFE7A3654850B5264D98833A10500041504C94679612B5A80612CC41956";
    attribute INIT_35 of inst : label is "C6989929C67510628C60BB9B924D580625D1596545A2618625DE3153A21683D8";
    attribute INIT_36 of inst : label is "DF9B61801773950784987194648112493D07021898699E50A991514326464289";
    attribute INIT_37 of inst : label is "B81464AA858696471419AA5A86A14722587092486E6966685B590F2E4DF5E003";
    attribute INIT_38 of inst : label is "A6422A4924940456208C2130C6458851D98414D3B1B9527884C485297185D334";
    attribute INIT_39 of inst : label is "8032892D0DFE219A00C1988855F908608E906162865F2228639988A2050A0A69";
    attribute INIT_3A of inst : label is "113D5D25F80317A5C5064F44DA40841133304116549BC71419A79907BBCA3554";
    attribute INIT_3B of inst : label is "985621E1281565993203E2569FFE00CA881F1882999886204593FE03641B9580";
    attribute INIT_3C of inst : label is "A88B0008988758A0A1DCAC664A6C5492958EB75E5A8BF9BFE2DC4D37C92F5488";
    attribute INIT_3D of inst : label is "99BAF38BC786A62908880D008262F0FA861099C0256265999FB028E662DA996D";
    attribute INIT_3E of inst : label is "BA26146B6649655410E4D34A81A8952106BC0444D18AC9C06E920944C00C3E88";
    attribute INIT_3F of inst : label is "E41AE60078B0780402C8266D6C6877E949DDC1150C8D1A7B30C3A9129B163658";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
