-- generated with romgen v3.0 by MikeJ
library ieee;
  use ieee.std_logic_1164.all;
  use ieee.std_logic_unsigned.all;
  use ieee.numeric_std.all;

library UNISIM;
  use UNISIM.Vcomponents.all;

entity GFX1 is
  port (
    CLK         : in    std_logic;
    ENA         : in    std_logic;
    ADDR        : in    std_logic_vector(13 downto 0);
    DATA        : out   std_logic_vector(7 downto 0)
    );
end;

architecture RTL of GFX1 is

  function romgen_str2bv (str : string) return bit_vector is
    variable result : bit_vector (str'length*4-1 downto 0);
  begin
    for i in 0 to str'length-1 loop
      case str(str'high-i) is
        when '0'       => result(i*4+3 downto i*4) := x"0";
        when '1'       => result(i*4+3 downto i*4) := x"1";
        when '2'       => result(i*4+3 downto i*4) := x"2";
        when '3'       => result(i*4+3 downto i*4) := x"3";
        when '4'       => result(i*4+3 downto i*4) := x"4";
        when '5'       => result(i*4+3 downto i*4) := x"5";
        when '6'       => result(i*4+3 downto i*4) := x"6";
        when '7'       => result(i*4+3 downto i*4) := x"7";
        when '8'       => result(i*4+3 downto i*4) := x"8";
        when '9'       => result(i*4+3 downto i*4) := x"9";
        when 'A'       => result(i*4+3 downto i*4) := x"A";
        when 'B'       => result(i*4+3 downto i*4) := x"B";
        when 'C'       => result(i*4+3 downto i*4) := x"C";
        when 'D'       => result(i*4+3 downto i*4) := x"D";
        when 'E'       => result(i*4+3 downto i*4) := x"E";
        when 'F'       => result(i*4+3 downto i*4) := x"F";
        when others    => null;
      end case;
    end loop;
    return result;
  end romgen_str2bv;

  attribute INIT_00 : string;
  attribute INIT_01 : string;
  attribute INIT_02 : string;
  attribute INIT_03 : string;
  attribute INIT_04 : string;
  attribute INIT_05 : string;
  attribute INIT_06 : string;
  attribute INIT_07 : string;
  attribute INIT_08 : string;
  attribute INIT_09 : string;
  attribute INIT_0A : string;
  attribute INIT_0B : string;
  attribute INIT_0C : string;
  attribute INIT_0D : string;
  attribute INIT_0E : string;
  attribute INIT_0F : string;
  attribute INIT_10 : string;
  attribute INIT_11 : string;
  attribute INIT_12 : string;
  attribute INIT_13 : string;
  attribute INIT_14 : string;
  attribute INIT_15 : string;
  attribute INIT_16 : string;
  attribute INIT_17 : string;
  attribute INIT_18 : string;
  attribute INIT_19 : string;
  attribute INIT_1A : string;
  attribute INIT_1B : string;
  attribute INIT_1C : string;
  attribute INIT_1D : string;
  attribute INIT_1E : string;
  attribute INIT_1F : string;
  attribute INIT_20 : string;
  attribute INIT_21 : string;
  attribute INIT_22 : string;
  attribute INIT_23 : string;
  attribute INIT_24 : string;
  attribute INIT_25 : string;
  attribute INIT_26 : string;
  attribute INIT_27 : string;
  attribute INIT_28 : string;
  attribute INIT_29 : string;
  attribute INIT_2A : string;
  attribute INIT_2B : string;
  attribute INIT_2C : string;
  attribute INIT_2D : string;
  attribute INIT_2E : string;
  attribute INIT_2F : string;
  attribute INIT_30 : string;
  attribute INIT_31 : string;
  attribute INIT_32 : string;
  attribute INIT_33 : string;
  attribute INIT_34 : string;
  attribute INIT_35 : string;
  attribute INIT_36 : string;
  attribute INIT_37 : string;
  attribute INIT_38 : string;
  attribute INIT_39 : string;
  attribute INIT_3A : string;
  attribute INIT_3B : string;
  attribute INIT_3C : string;
  attribute INIT_3D : string;
  attribute INIT_3E : string;
  attribute INIT_3F : string;

  component RAMB16_S1
    --pragma translate_off
    generic (
      INIT_00 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_01 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_02 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_03 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_04 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_05 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_06 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_07 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_08 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_09 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_0F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_10 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_11 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_12 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_13 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_14 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_15 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_16 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_17 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_18 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_19 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_1F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_20 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_21 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_22 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_23 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_24 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_25 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_26 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_27 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_28 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_29 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_2F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_30 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_31 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_32 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_33 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_34 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_35 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_36 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_37 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_38 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_39 : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3A : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3B : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3C : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3D : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3E : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000";
      INIT_3F : bit_vector (255 downto 0) := x"0000000000000000000000000000000000000000000000000000000000000000"
      );
    --pragma translate_on
    port (
      DO    : out std_logic_vector (0 downto 0);
      ADDR  : in  std_logic_vector (13 downto 0);
      CLK   : in  std_logic;
      DI    : in  std_logic_vector (0 downto 0);
      EN    : in  std_logic;
      SSR   : in  std_logic;
      WE    : in  std_logic 
      );
  end component;

  signal rom_addr : std_logic_vector(13 downto 0);

begin

  p_addr : process(ADDR)
  begin
     rom_addr <= (others => '0');
     rom_addr(13 downto 0) <= ADDR;
  end process;

  rom0 : if true generate
    attribute INIT_00 of inst : label is "784088773F3CFF0020A0403B2F23001101980007007400F7FF000000FF000000";
    attribute INIT_01 of inst : label is "1FFEF03F1FE1F00F05FE401F050140004410613CAA0A5550AA2A555455555555";
    attribute INIT_02 of inst : label is "FC00440000D10000F89F030700E20078F998030700C400F100008A04FE440000";
    attribute INIT_03 of inst : label is "3C00100030304800002000183F003C000C007E00030066001E001E000C006300";
    attribute INIT_04 of inst : label is "63007F007F003000780003000C007F0067007E003E00630060007E006300A13C";
    attribute INIT_05 of inst : label is "000000000000000000181C001E001C007F00770063000C003E00670063006300";
    attribute INIT_06 of inst : label is "4438C66B36BC16C86E00D200B65CCAF27E00FB00F65EEAF27E00FF00FE5EFBF2";
    attribute INIT_07 of inst : label is "00B300650000000048A22430000000001838195B00400004C2BA92BB68DA531D";
    attribute INIT_08 of inst : label is "1000100000000020200011000848177A000000000040071A0000000000000618";
    attribute INIT_09 of inst : label is "0000000000000000C60038000029004500F802FF8080FFFFFEF8FFFF038000FF";
    attribute INIT_0A of inst : label is "2000010100070087004010101C42000080700902004002000000800083008780";
    attribute INIT_0B of inst : label is "00030202C8020300000003080000844EC000636000C400930001208000000700";
    attribute INIT_0C of inst : label is "585810688C0088A40810010120600400202022009C80000096080300040000FF";
    attribute INIT_0D of inst : label is "9E8F08C0E0001101806000044090104818000000CCAF274E01024C27000320BC";
    attribute INIT_0E of inst : label is "44386000000F0200080010000000000080800B09CF0000E02E0F02E093010002";
    attribute INIT_0F of inst : label is "34FB6CB162D90D36ECECD9CFFCFCCFD9F8FCDFCFFCF8CFDFECCC3FFFFCF0CFDF";
    attribute INIT_10 of inst : label is "0F400C00F80348781FC0121EF0023000004406000003007C00C40C3E00020000";
    attribute INIT_11 of inst : label is "006C061F0003007C1E402C003C0102000F1803071C3820F01F0006187138000E";
    attribute INIT_12 of inst : label is "671F630788C0007807FFC60099C0003C1FC01E00F006F0000F49003FF8C90080";
    attribute INIT_13 of inst : label is "0000000000000000380000000000000000000000000000000000190000009800";
    attribute INIT_14 of inst : label is "0000000000000000000C06000000000000302000000000000000060000000000";
    attribute INIT_15 of inst : label is "0013000000000000000606000000000000380000001C0000000D0C0000B03000";
    attribute INIT_16 of inst : label is "001904001FF100000001C8E000F6001800000000080000001000000000000200";
    attribute INIT_17 of inst : label is "0000403C000602780060401E0000023CF00FF03F1FE11FFE4000403F050105FE";
    attribute INIT_18 of inst : label is "6F61000022550000E64E00002255000008490000C62900001C090000C6290000";
    attribute INIT_19 of inst : label is "C080000000011F000080F80003010000311C0207F8F008F061E5000022550000";
    attribute INIT_1A of inst : label is "C0E000000000000007000000B040000000D8000006C0001E6003067800933000";
    attribute INIT_1B of inst : label is "0001001F0080300000010C00008800F800040C000000003C0008183C00000000";
    attribute INIT_1C of inst : label is "0007000000E00000000E00000070000000040C07000000E0800E00180500001C";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000010000008000000003000000C00000";
    attribute INIT_1E of inst : label is "120000E7900000CE000000D200000096FF000000FE0000008140021FEC2300CF";
    attribute INIT_1F of inst : label is "07800E1EE001F0780FE100F0F0C7000F0F330E00E0C0E01001010000E6E71C10";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF00F87EFF000FF0FF07FFFFFFFFFF0000FFFFFFFF";
    attribute INIT_21 of inst : label is "00FF0CFF000F00FFE0FFFFFFFFFFFFFFFFFFFFFF3FFF00FF00FF003F00FFFEFF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF003F0000";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFF00FF00FFFFFFFFFFFFFFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF7FFFF800FFFFFFFF03FF00FF0000F880FFFF3FFF003FF0C0FFFFFFFF";
    attribute INIT_28 of inst : label is "FF00FF003F0000000000FF00FFC0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF07C000";
    attribute INIT_29 of inst : label is "FFFFFFFFE0F0FFFF00E0F0FFFFFF00FC00FFFFFFFFFFC0FEFFFFFF00FF00FF00";
    attribute INIT_2A of inst : label is "FFFFFFFFF000FFFFFFFFFFFFFFFFFFFFFFFF03FFC0FF00FFF0FFFFFF00F8FCFF";
    attribute INIT_2B of inst : label is "FFFF0701C000FFFFFFFFFFFF7F1FFCF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FF000300FFFFFFFFFFFFFFFFF8F8FFFFFFFFFFFFFFFF1F01FCF8FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFF0FFF000F000000FCFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F0080FFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "00200000000300000040000000040000004003000003307800C00C1E0002C000";
    attribute INIT_31 of inst : label is "0009000070C800000E130000009000000021000000C200000043000000840000";
    attribute INIT_32 of inst : label is "00040000002000000000000000000000030400006010000006080000C0200000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000020000004000000002000000400000";
    attribute INIT_34 of inst : label is "00200000000300000040000000040000004000000003007C00C0003E00020000";
    attribute INIT_35 of inst : label is "00080000700800000E1000000010000000200000000200000040000000040000";
    attribute INIT_36 of inst : label is "0000000018300000200000006230000000000C071C3820F0000000187138000E";
    attribute INIT_37 of inst : label is "01000000806000000C1000005860000000000000906000001000000054600000";
    attribute INIT_38 of inst : label is "0006000000600000000100000080000000060000006000000001000000800000";
    attribute INIT_39 of inst : label is "0000000000000000000000000000000000060000006000000001000000800000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "00060000000000000000000000000000000C0000000000000000000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(0 downto 0),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom1 : if true generate
    attribute INIT_00 of inst : label is "704022143F3CFF002020400A213D001B009C000000700087FFFF0000FFFF0000";
    attribute INIT_01 of inst : label is "EFFFEF7E3FE3F88F0103000004016040929201065555AAAA54552AAAAAAAAAAA";
    attribute INIT_02 of inst : label is "FD06490400800004F898030000080042F89C0300001000840000F28AFE6C0000";
    attribute INIT_03 of inst : label is "0000080030306C0000100018633C723E0618603E7E3E36060C3E077F0C3F631C";
    attribute INIT_04 of inst : label is "633E7B637F63303F6C67033E0C3F6363601F6060303F637C601E637E63639D42";
    attribute INIT_05 of inst : label is "FF006100FD003F0000180E7F330C3E636B636308633E0C0C603E6367633D6360";
    attribute INIT_06 of inst : label is "31929A1A52C9D11DE4BCCE7B76BA37EDEEFCEE7F7EBAB7FDFEFCFE7FFEBEF7FD";
    attribute INIT_07 of inst : label is "00040021000000004008008400000000C64D45960000000008B00C99508106D4";
    attribute INIT_08 of inst : label is "140028000004001014400A008044001100000000804000110000000000000018";
    attribute INIT_09 of inst : label is "FC003F00F000FF00290045000029007900F0027F8080FFFFFEF8FFFF038000FF";
    attribute INIT_0A of inst : label is "3000010100F80080003020100081000000F01004004004000000700000007880";
    attribute INIT_0B of inst : label is "0004010290023F008000E104000003270300187E00020008001E207C80000700";
    attribute INIT_0C of inst : label is "98580830820E84A40410010120700400102021009C80000027080F0002C00000";
    attribute INIT_0D of inst : label is "9E8F0420C0001302800000025080082006000007CCAE274E01024CCE0000405C";
    attribute INIT_0E of inst : label is "319210000070040004C0200300000000808009CB9E1F001C2C10011093020001";
    attribute INIT_0F of inst : label is "6CFA6CD9C2D20616ECECD9DF0000E0D8F8FCDFDF0000E0D8CCEC7FFF0000E0D8";
    attribute INIT_10 of inst : label is "0FC3061CF8E1307C1F470C3EF0C4603800C6031C0001007C004C063E00040038";
    attribute INIT_11 of inst : label is "006C0000000300001C4000001C0100001F0006031C3800E01FEE003878380046";
    attribute INIT_12 of inst : label is "7F100F0100C000980EB106000080000C9F470C00F2C460F80769003FF04B00BC";
    attribute INIT_13 of inst : label is "0000003000000000000000000000000000000000000000000000180000001800";
    attribute INIT_14 of inst : label is "181C000000000000000C03000000000000302000000000000004040000800000";
    attribute INIT_15 of inst : label is "00020000000000000063000000000000001C0000003800000019000000980000";
    attribute INIT_16 of inst : label is "180100031BE000F81C01043C18EC001C042000004C0400003200000020000000";
    attribute INIT_17 of inst : label is "001846180006006000680C0600000218EF8FF87EEFE33FFF0040600001010503";
    attribute INIT_18 of inst : label is "9811000055550000494800005555000009290000292900000909000029290000";
    attribute INIT_19 of inst : label is "C606000000033F0018CCFC0003000000311C0303F800B8E09185000055550000";
    attribute INIT_1A of inst : label is "E0C300000080000007040000B0400000401E000002F0001E4003007802180000";
    attribute INIT_1B of inst : label is "0011001F0090000000080000004800F8000C06000000003800180C1C00000000";
    attribute INIT_1C of inst : label is "0007000000E00000000E000000700000000E0001000000C00046003800000006";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000003000000C00000";
    attribute INIT_1E of inst : label is "120000C0900000060000000C000000607F000000FC0000008100000FC01848FC";
    attribute INIT_1F of inst : label is "8FE7060CF1C7603007890060E04100061F010603E88040F800010000FCC20C18";
    attribute INIT_20 of inst : label is "7FFFF0FFFFFFFFFFFFFFFF0000E018FF0007C0FE037F0000FFFF0000FFFFFFFF";
    attribute INIT_21 of inst : label is "00F800FF000300FC80FFFFFFFFFFFFFFFEFFFFFF0FFF00FF00FF000C00F8F8FF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFF001F0000";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFDFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFF00FFFFFFFFFFFFFFFFFFFFFF0FFFFCFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF3FFFFC00FFFFFFFF00FF003F0000FEE0FFFF0FFF000FF0F0FFFFFFFF";
    attribute INIT_28 of inst : label is "FF00FF00FF000000C000FF00FFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FE000";
    attribute INIT_29 of inst : label is "FFFFFFFFE0F0FFFF00C080FFFFFF00F000FF00FFFFFF00FEFFFFFFFFFF00FF00";
    attribute INIT_2A of inst : label is "FFFF07010000FEFCFFFFFFFFFFFF7F1FFFFF033F80FE00FC00FFFFFF00C0FFFF";
    attribute INIT_2B of inst : label is "3F0300000000FFFFFFFFFFFF00000000F8F8FFFFFFFFFFFFFFFFF8F8FFFFFFFF";
    attribute INIT_2C of inst : label is "000000000080FFFFFF0701000000FCFEFFFFFF7F1F0000000000FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FEFFFFFFFFFF00000000000000000000F0F8FFFFFFFFC0E0FFFFFFFFFF0F0F00";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000000080";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0061000000E100700007000E0080000000C3001C00E1007C0047003E00C40038";
    attribute INIT_31 of inst : label is "001100000044000000020000008000000032000000A600000025000000480000";
    attribute INIT_32 of inst : label is "00000000C0000000030000000000000000080000600800000600000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "00600000000100780000001E0000000000C0001C0001007C0040003E00040038";
    attribute INIT_35 of inst : label is "0010000000040000000000000000000000300000000600000020000000080000";
    attribute INIT_36 of inst : label is "00000003187000F0003600087030000C000000031C3800E000E0003878380046";
    attribute INIT_37 of inst : label is "0000000010600000080A00006840000000000000106000000018000064600000";
    attribute INIT_38 of inst : label is "00000000000000000007000000E0000000000000000000000007000000E00000";
    attribute INIT_39 of inst : label is "0000000000000000000100000080000000000000000000000005000000A00000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "00000000000000000036000000000000000C000000000000006C000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000000000000000000000000000000000018000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(1 downto 1),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom2 : if true generate
    attribute INIT_00 of inst : label is "604036803C3F3CFF6020440A3F3D001B8226000100700007FFFF0000FFFF0000";
    attribute INIT_01 of inst : label is "E77FCFFC7EE7FCCF013900301801304010443003AAAA5555AA2A555455555555";
    attribute INIT_02 of inst : label is "FF7F491E00080003F220010100080002F22601010010000400000492387C0000";
    attribute INIT_03 of inst : label is "00000C0030006C0000300000630662436318306360631E06066363701C0C2632";
    attribute INIT_04 of inst : label is "6363736777633030666E03630C0C63633033606030306666333363633663429D";
    attribute INIT_05 of inst : label is "FF00B100FD007F0000000770330C77776377631C63630C0C6663636E63666360";
    attribute INIT_06 of inst : label is "E2A20C9968DA63DDF2D2BEBB72DAF7DDF2DABEFB7ADEF7FDF2DEBEFBFEDEF7FD";
    attribute INIT_07 of inst : label is "000000000000000000200011000000001020904200000000B44C644A00360086";
    attribute INIT_08 of inst : label is "0A0060000008003888800C000048011A00000C000050011A0000080000000000";
    attribute INIT_09 of inst : label is "FC007F00F800FF002900050000290041000002028080FFFF00FC00FF0001007F";
    attribute INIT_0A of inst : label is "3000020100000000000F20100081000000E020040080380000000F0000000080";
    attribute INIT_0B of inst : label is "0000010220041E00E0007004E0C00033FC00073F0003000700E02043C0000100";
    attribute INIT_0C of inst : label is "18580810420F84900408010140B00201102011009C98800027881C0002300000";
    attribute INIT_0D of inst : label is "9E9F041080602304A01800015080082001C00000CCCE234E0102444E00008020";
    attribute INIT_0E of inst : label is "E2A208000080040004204004F0000F00C080093B9C200002CC23000897040001";
    attribute INIT_0F of inst : label is "68362CD8C1B2071B0C6CD8D8FC007FD80000C0D8FC007FD81C6CE000FC007FD8";
    attribute INIT_10 of inst : label is "078F0003F0F900FC8F1F003FE1F000C0008600000001007C800C003E01000000";
    attribute INIT_11 of inst : label is "00400000000100000060061E0003003C1F6600001C7000441E63006738300063";
    attribute INIT_12 of inst : label is "3E000600000000CC7E000C00000000C68F53003CE29400F8034F003FE07900F0";
    attribute INIT_13 of inst : label is "00000030000000001800000000000000000033000000CC0000000C0000003000";
    attribute INIT_14 of inst : label is "380E000000000000000C00000000000000000000000000000004000000800000";
    attribute INIT_15 of inst : label is "4E00000000000000002300000000000001000000800000000018000000180000";
    attribute INIT_16 of inst : label is "300CC0077B0000FD3C0C001F781800060C000000380000001C00000030002000";
    attribute INIT_17 of inst : label is "004C420808020080104C060100020210CFCFFCFCE7E77E7F0040303001011839";
    attribute INIT_18 of inst : label is "149900005555000049C90000555500007D190000292900000919000029290000";
    attribute INIT_19 of inst : label is "CE03000000023F003846FC0003000000390C0111F8F090009F930000D5550000";
    attribute INIT_1A of inst : label is "FF11000080800000030D000320C00040C11E000082F0000E400F007003780000";
    attribute INIT_1B of inst : label is "001E000E001800340018002C00780070000C000C000000380018001C00000030";
    attribute INIT_1C of inst : label is "00020000004000000006000000600000004600000000004000C6006400000002";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0C000047600000C400000000000000000F00001CE0000070C0000083980000F8";
    attribute INIT_1F of inst : label is "8FE30004F197002000890047004100E23D080007D02000E8000000007810001E";
    attribute INIT_20 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFF00C000FF000380FC013FFFFFFFFF0000FFFFFFFF";
    attribute INIT_21 of inst : label is "00C000FF000000F000FFFFFFFFFF7FFFF0FFFFFF07FF000300FF000000E0E0FF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF070300";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF1FFFFEC0FFFF0FFF00FF000FC000FFF0FFFF03FF0003F0F0FFFFFFFF";
    attribute INIT_28 of inst : label is "FFFFFF0FFF000F00F000FF00FFFCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF7FF080";
    attribute INIT_29 of inst : label is "FFFFFFFFE0F0FFFF008000FFF8FF000000FF00FFFFFF00FEFFFFFFFFFF00FFF0";
    attribute INIT_2A of inst : label is "FFFFFFFFFCC0FFFFFFFFFFFFFFFFFFFF9FFF010F00FC00E000FFF0FFC000FFF0";
    attribute INIT_2B of inst : label is "FFFF0F03E080FFFFFFFFFFFFFF3FFEF8FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2C of inst : label is "FF3F3F00FFFFFFFFFFFFFFFFF8F8FFFFFFFFFFFFFFFF7F07FEF8FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FFFFFFFFFFFFFFFFFF0FFF000F00F8FCFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0080FEFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "0043000E00F10078800F001E02C000700081000000C1007C8003003E01800000";
    attribute INIT_31 of inst : label is "000000000000000000000000000000000023000E006200784006001E04C00070";
    attribute INIT_32 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000800000000100000000000000";
    attribute INIT_34 of inst : label is "0040000E000100788000001E02000070008000000001007C8000003E01000000";
    attribute INIT_35 of inst : label is "000000000000000000000000000000000020000E000200784000001E04000070";
    attribute INIT_36 of inst : label is "00160001386000E00016001870200044006000001C700044006C006438300063";
    attribute INIT_37 of inst : label is "001A000030400000000000006000000000080003306000C0000A000C60400018";
    attribute INIT_38 of inst : label is "0100000080000000000600000060000001000000800000000006000000600000";
    attribute INIT_39 of inst : label is "0100000080000000000200000040000001000000800000000006000000600000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "200000000000000000160000000000004000000000000000002C000000000000";
    attribute INIT_3F of inst : label is "0000000000000000000D0000000000001000000000000000000B000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(2 downto 2),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom3 : if true generate
    attribute INIT_00 of inst : label is "40C000803C3F3CFF7F204440002300008203700000200003FFFF0000FFFF0000";
    attribute INIT_01 of inst : label is "E33F8FF8FCEF7EEF010D0040000100400000006150550AAA54552AAAAAAAAAAA";
    attribute INIT_02 of inst : label is "F9F9093000300000F2F0390100B00001E2F3730100200003F800F8FA107C0000";
    attribute INIT_03 of inst : label is "003C0C0030306C00003000003E033C4F7F181E637E030E7F3F033E3C0C0C1C63";
    attribute INIT_04 of inst : label is "3E63636F636B3030637C03033F0C63631F637F603F307C631E607E631C7F3CA1";
    attribute INIT_05 of inst : label is "0100B0000D00E00000007F38330C633E637F633E63633F0C3C037E7C3E6F7E7E";
    attribute INIT_06 of inst : label is "086C64C270830640EEAE4EBDFCCA6EDDEEBECEBDFCDE7FDDEEBECEFDFCDE7FFD";
    attribute INIT_07 of inst : label is "00000000000000000009004100000000648A43C4000000004931C9D6005200D4";
    attribute INIT_08 of inst : label is "0408700800000010B0801C0200B0000E20001C0000A0000E000018000000000C";
    attribute INIT_09 of inst : label is "0000E0001C0000002900050000C6007C000002028080FFFF00FC00FF00010000";
    attribute INIT_0A of inst : label is "7000020100000000000020100062000000C040090000C001FF000000007C0080";
    attribute INIT_0B of inst : label is "00000102C0C400009800B8061FE0004800F0008F00FC000000001020C0003C00";
    attribute INIT_0C of inst : label is "305808103C738290040802018040010208200E1C4C98C0006790000101080000";
    attribute INIT_0D of inst : label is "9E9E020800E02708B0E000005040881000200000CCCE114E0101404E0000801E";
    attribute INIT_0E of inst : label is "086C048080000901021040080F00F000C080040B984F00014C270004A7090001";
    attribute INIT_0F of inst : label is "5834345880A2030BFC6CD9D8FCFC3FDFF800DFD8FCFC3FDFF86CCF00FCFC3FDF";
    attribute INIT_10 of inst : label is "430C0007E14800F08712000FC33000E040000000010000008000000003000000";
    attribute INIT_11 of inst : label is "484C000001010000402C001E0102003C1EE300073870000C1803004F38200075";
    attribute INIT_12 of inst : label is "1F2300438000008EFF5E0003800000CF8712000FC29000E04346000FE13100F8";
    attribute INIT_13 of inst : label is "00000000000000000C0000180000000000000000000000000001000000800000";
    attribute INIT_14 of inst : label is "3800000000000000000000000000000000200000000000000004000000000000";
    attribute INIT_15 of inst : label is "DF00000000000000000F000000000000390000009C000000001E000000780000";
    attribute INIT_16 of inst : label is "302C0C0FF3000003240C300FF7000083070200000020000000800800E0000000";
    attribute INIT_17 of inst : label is "006000100C020000304C0000000600088FEF7EF8E3EFFC3F004000400101000D";
    attribute INIT_18 of inst : label is "126600005522000049460000552200004908000029C600000908000029C60000";
    attribute INIT_19 of inst : label is "8E0000C001061E00B86078000100000339060031F86800F09961000055220000";
    attribute INIT_1A of inst : label is "FF310000C080000000000007808000E0C90C0000C0600004410F002083780000";
    attribute INIT_1B of inst : label is "000C000400780024011E00248030002000000000000000180000001800000000";
    attribute INIT_1C of inst : label is "00000000000000000D000000B000000000C6000000000000040C00C000000003";
    attribute INIT_1D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_1E of inst : label is "0000005F000000F400000000000000000300007E800000FC40000080220100F8";
    attribute INIT_1F of inst : label is "87020004E1900020E386006FE76100F638080007102000E800000001F81000E0";
    attribute INIT_20 of inst : label is "07FFE0FFFFFFFFFFFFFFFFFF008000FF000000F8001F0000FFFF0000FFFFFFFF";
    attribute INIT_21 of inst : label is "0000003E0000000000FCFCFFFFFF1FFFC0FFFFFF03FF000000000000008000FF";
    attribute INIT_22 of inst : label is "FFFFFFFFFFFFFFFF80FFFFFFF0FFFFFFFFFFFFFFFFFFFFFFFFFF0FFF00010000";
    attribute INIT_23 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF3FFFE0FFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_25 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_26 of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_27 of inst : label is "FFFFFFFF03FFFFF0FFFF00FF001F0000FC00FFF0FFFF00FF0000F0F0FFFFFFFF";
    attribute INIT_28 of inst : label is "FFFFFFFFFF07FF00FC00FF00FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFCC0";
    attribute INIT_29 of inst : label is "FFFFFFFFE0F0FFFF000000FEC0FF000000FF00FFFFFFF0F0FFFFFFFFFFFFFFFF";
    attribute INIT_2A of inst : label is "FFFF0F030000FEFCFFFFFFFFFFFFFF3F00FF000700F0000000FC00FFE000FFF8";
    attribute INIT_2B of inst : label is "FF0F00000000FFFFFFFFFFFF00000000F8F8FFFFFFFFFFFFFFFFFCF8FFFFFFFF";
    attribute INIT_2C of inst : label is "000000000080FFFFFF3F0F000000FCFEFFFFFFFFFF0300000000FFFFFFFFFFFF";
    attribute INIT_2D of inst : label is "FCFFFFFFFFFF00000000000000000000F0F8FFFFFFFFC0E0FFFFFFFFFFFFFF00";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00FF0000000000";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "2003000002300078C00C001E06C000004003000001300000800C000003C00000";
    attribute INIT_31 of inst : label is "00000006000000702000000E0800006000000000000000784000001E04000000";
    attribute INIT_32 of inst : label is "0000000000000000040000002000000000000000000000001000000010000000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "2000000002000078C000001E0600000040000000010000008000000003000000";
    attribute INIT_35 of inst : label is "00000006000000702000000E0800006000000000000000784000001E04000000";
    attribute INIT_36 of inst : label is "0036000038600048000000343000006A00EC00003870000C000C004038200075";
    attribute INIT_37 of inst : label is "00000003300000C00000000660000030001A0001304000800000001C60000048";
    attribute INIT_38 of inst : label is "07000000E0000000000000000000000007000000E00000000000000000000000";
    attribute INIT_39 of inst : label is "0200000040000000000000000000000005000000A00000000000000000000000";
    attribute INIT_3A of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3C of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3D of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_3E of inst : label is "66000000000000000000000000000000C0000000000000000000000000000000";
    attribute INIT_3F of inst : label is "1A00000000000000000000000000000036000000000000000000000000000000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(3 downto 3),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom4 : if true generate
    attribute INIT_00 of inst : label is "0000FF770000000080807F3B00801F35FD980707F09C07FCFF00FF0000000000";
    attribute INIT_01 of inst : label is "FE00FF00FE1EFFF0FE00FF20FEFEFFFF4410FE00FF0EFF70FE3E7F7C7F7FFFFF";
    attribute INIT_02 of inst : label is "FC001F00003C073CFC000700F81C0307FC000700F038070E00000000FE440000";
    attribute INIT_03 of inst : label is "3C00100030304800002000183F003C000C007E00030066001E001E000C006300";
    attribute INIT_04 of inst : label is "63007F007F003000780003000C007F0067007E003E00630060007E006300A13C";
    attribute INIT_05 of inst : label is "000000000000000000181C001E001C007F00770063000C003E00670063006300";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "2E006E001C1F38DCDC002E00F0B60A1DFC003F00F8BE1A7DFC003F00F8FE1F7F";
    attribute INIT_09 of inst : label is "0000000000000000C600380000290045F0F87FFF8080FFFF00000000008000FF";
    attribute INIT_0A of inst : label is "FFFF000000F80000003FE0E0E381FFFFFFFF07010080FCFFFFFF7FFF00FF787F";
    attribute INIT_0B of inst : label is "FFFC0101F0FCFFFFFFFFFCF7FFFF03BFFFFF1FFF00FB000F00FEC07FFFFFFFFF";
    attribute INIT_0C of inst : label is "BFBFEF9703FF071F070FFEFE1FFFF8FFDFDFC1FF7F7FFFFFEFF7FFFFFBFFFF00";
    attribute INIT_0D of inst : label is "7F7FF000FFFFEFFE7FFFFFFBBF7FEFBFE7FFFFFF3F1F1F3FFEFCBFDFFFFCDF7F";
    attribute INIT_0E of inst : label is "00008000FF000100F0000F0000000000FFFFF7073F00FF001F00FC000F00FFFC";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "3F3F1C00FEFCCC007F3F3300FCFC38003F3F1F00FEFCFC007F3F3F00FCFCF800";
    attribute INIT_11 of inst : label is "3F1F0F00FEFCF800013F1F00C0FEFC000F1F1300E2C4DC001F1F1F008CC4FC00";
    attribute INIT_12 of inst : label is "07181300F43EF80007002700E03EF0003F3F3F00F8F8F8003F381F00FE0EFC00";
    attribute INIT_13 of inst : label is "0000007F000000FEFF1F001FFFF800F800007F000000FE00007FF80000FE1F00";
    attribute INIT_14 of inst : label is "FF7F073FFFFEE0FC3F7F3F00FCFEFC00F0E0F06000000000FFFF7F1E80808000";
    attribute INIT_15 of inst : label is "7F33031FFFFEE0FC1F3F1F00FCFEF800FF79073FFF9EE0FC3F7E3F00FC7EFC00";
    attribute INIT_16 of inst : label is "FF7F003FE0F000F8FF67C01FF8F000E0FF07007FCFF000FEF30F007FFFE002FE";
    attribute INIT_17 of inst : label is "7FFF1F00E0F8F800071F1F00FEFFF800FFF0FF00FE1EFE00FFFFFF00FEFEFE00";
    attribute INIT_18 of inst : label is "6F61000022550000E64E00002255000008490000C62900001C090000C6290000";
    attribute INIT_19 of inst : label is "FF7F0F0FFFFFCCFCFFFF3300FFFEF8000E231E00FCFC4C0061E5000022550000";
    attribute INIT_1A of inst : label is "0F0F0F00FEFFFE00000200007F7FFCFE3F393F00FECEFC0067723F00F81CFC00";
    attribute INIT_1B of inst : label is "5F723F1FF57FFE00AFFE7F00FA4EFCF82F7F3F00FBFFFE3CDFFF7F3CF4FEFC00";
    attribute INIT_1C of inst : label is "0F1F0300F0F8C0001F3F0F00F8FCF0003F7F3F07EAFEFCE0BF7F3F18F5FEFC1C";
    attribute INIT_1D of inst : label is "00010000008000000003000000C000000007000000E00000030F0000C0F00000";
    attribute INIT_1E of inst : label is "3307001F98C000F00000003300000098FF000000FE0000003E3F021F1CE400C0";
    attribute INIT_1F of inst : label is "1F3F1F00F8FCF8003F1E0F00FC38F000F04C7F00E030F000FF3E0F00E018FF00";
    attribute INIT_20 of inst : label is "F787011FFFFFC31F03000000FFFF9FFFFFF1FFFFF9030000FFFFFFFF0000FFFF";
    attribute INIT_21 of inst : label is "FFFFFF1FFFF0FFFFFFFFFFF7DFFF0000FEC00F3FC0FFFFFFFFFFFFC7FFFFFFFF";
    attribute INIT_22 of inst : label is "FFF0FFFF7FFFE0FFFFFFFFFFF07F01F807FF0FFF60FFFFFFF8C70710FFC0FFFF";
    attribute INIT_23 of inst : label is "00FF01FFFFFF2FFFF1FFBFFF83FF3FFF00FFFFFF7FFF00FFFFFF8F1F0300E100";
    attribute INIT_24 of inst : label is "FF0FFF00FF00FF00FFFCFFFF07FFC0FFFFFFFFFFFF1FFF0000FE00FFFFFF00FF";
    attribute INIT_25 of inst : label is "F0FFFFFFFFFFFFFF0FFF00FFFFFFFFC3FF00FFFF3FFF00FFE0FFFF00FFFCFF00";
    attribute INIT_26 of inst : label is "00FF00FF00FF00FF00FF00000000FF000FFF00FF00FFFFFFFFFFFF00FF00F3DF";
    attribute INIT_27 of inst : label is "C000F800FF7F07FFC000FFFFFFFFFFFFFFFF077FFC00FFFFFFFF0F3FFF0000FF";
    attribute INIT_28 of inst : label is "00FF00FFC0FFFFFFFFFF00FF003FC000FFF80F00F8001F000000000000F83FFF";
    attribute INIT_29 of inst : label is "00FF00FF1F0FFFF0FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFE1FFFF00FF00FF00FF";
    attribute INIT_2A of inst : label is "3F0F00000FFF0000E0E0FFFF7F3F0000FFFFFFFFFFFFFFFFFFFFFFFFFFFF03FF";
    attribute INIT_2B of inst : label is "0000F8FE3FFFF8FEFFFF1F0180E0030F0000E0F0FFFFFFFF03010000FFFFFFFF";
    attribute INIT_2C of inst : label is "00FFFCFF0000FFFF0000000007070000FFFF00000000E0FE030780E0FFFFFFFF";
    attribute INIT_2D of inst : label is "0000FFFFFF0300F000FFF0FFFFFF03010000FFFFFFFF0000FF03030000000000";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00E0F8000000F0FF7F0000";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "1F1F1900FCFCCC003F3F3300F8F898003F3F1300FEFCB4007F3F2D00FCFCC800";
    attribute INIT_31 of inst : label is "070603008030E000010C0700E060C0001F1E0700FC3CF0003F3C0F00F878E000";
    attribute INIT_32 of inst : label is "0002000000C000000002000000C000000002000000E000000005000000C00000";
    attribute INIT_33 of inst : label is "0000000000800000000100000000000000010000008000000001000000800000";
    attribute INIT_34 of inst : label is "1F191C00FCFCFC003F333900F8F8F8003F3B1900FEFCFC007F3B3300FCFCF800";
    attribute INIT_35 of inst : label is "0705030080F0E000010B0700E0E0C0001F1C0700FCFCF0003F390F00F8F8E000";
    attribute INIT_36 of inst : label is "030F0900E0C8F800070F070098C8F0000F1F1C00E2C4DC001F1F19008CC4FC00";
    attribute INIT_37 of inst : label is "000703000090E00003040000A0900000000707000090F00003070300A090E000";
    attribute INIT_38 of inst : label is "7F270000FEE400001F3A1B00F85CD800FF47073FFFE2E0FC3F723300FC4ECC00";
    attribute INIT_39 of inst : label is "1F090000F8900000000F030000F0C0003F170000FCE80000071E0F00E078F000";
    attribute INIT_3A of inst : label is "00000000000000000003000000C0000007070000E0E000000007000000E00000";
    attribute INIT_3B of inst : label is "0000000000000000000100000000000000010000008000000003000000800000";
    attribute INIT_3C of inst : label is "7F230000FEFC00001F391C00F8FCF800FF7F073FFFFEE0FC3F733900FCFEFC00";
    attribute INIT_3D of inst : label is "1F0D0000F8F00000000D030000F0C0003F190000FCF80000071D0F00E0F8F000";
    attribute INIT_3E of inst : label is "3F1E0000FEFC0000071C0F00F0FCF8007F2C031FFFFEE0FC1F391900FCFEF800";
    attribute INIT_3F of inst : label is "0F070000F8F000000007010000F0C0001F0F0000FCF80000030F0300E0F8F000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(4 downto 4),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom5 : if true generate
    attribute INIT_00 of inst : label is "00006B140000000080007F0A0080003FFC9C0700E098038CFFFFFFFF00000000";
    attribute INIT_01 of inst : label is "1EFCF07FFE1EFFF0FEFCFF7FFFFEFFFF9292FE78FF7FFFFEFE7F7FFEFFFFFFFF";
    attribute INIT_02 of inst : label is "FCE0380000F8001CFC000700F04C0106FC000700E098030C00000000FE6C0000";
    attribute INIT_03 of inst : label is "0000080030306C0000100018633C723E0618603E7E3E36060C3E077F0C3F631C";
    attribute INIT_04 of inst : label is "633E7B637F63303F6C67033E0C3F6363601F6060303F637C601E637E63639D42";
    attribute INIT_05 of inst : label is "000000000000000000180E7F330C3E636B636308633E0C0C603E6367633D6360";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "6BF0B50F101B08AAE880350370BA0F6EFCC03F0370BE0F6EFCC03F03F0FE0F7F";
    attribute INIT_09 of inst : label is "00000000000000002900450000290079F0F07F7F8080FFFF00000000008000FF";
    attribute INIT_0A of inst : label is "FFFF000000000000000FC0E0FF00FFFFFFFF0F030080F8FFFFFF0FFF00FF007F";
    attribute INIT_0B of inst : label is "FFFB0001E0FCFFFF7FFFFEFBFFFF00DFFCFF07FF00FD000700E0C083FFFFFFFF";
    attribute INIT_0C of inst : label is "7FBFF7CF01FF031F030FFEFE1FFFF8FFEFDFC0FF7F7FFFFFDFF7FFFFFD3FFFFF";
    attribute INIT_0D of inst : label is "7F7FF8C0FFFFEFFD7FFFFFFDBF7FF7DFF9FFFFF83F1F1F3FFEFCBF3FFFFFBFBF";
    attribute INIT_0E of inst : label is "0000E000FF0F0300F8001F0000000000FFFFF7077F00FFE01F0FFEE00F01FFFE";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "3F1C1F00FE1CFC007F383F00FC38F8003F1F1F00FEFCFC007F3F3F00FCF8F800";
    attribute INIT_11 of inst : label is "3F1F030FFEFCE0F8033F3F00E0FEFE001F1F1F00E2C4FC001F1F0F0086C4F800";
    attribute INIT_12 of inst : label is "071F1F00FE3CF8000F3E2700FC7EF0007F383F00FC38F8003F190F00FECCF800";
    attribute INIT_13 of inst : label is "000000FF000000FFFF00007FFF0000FE0000FF000000FF0000FFF90000FF9F00";
    attribute INIT_14 of inst : label is "FF7F007FFFFE00FE3F7F1F00FCFEF800F0E0F0F000000000FFFF7F3F80000000";
    attribute INIT_15 of inst : label is "7F13003FFFFE00FE1F130F00FCFEF800FF7F007FFFFE00FE3F781F00FC1EF800";
    attribute INIT_16 of inst : label is "FF3F007CF8E00000FF3F0443F8E000E07C2000FFCF0400FFF30000FF3E0000FF";
    attribute INIT_17 of inst : label is "FF7F1F00E0F8F800071F1F00FFFEF800F0F0FF7F1E1EFEFCFFFFFF7FFEFEFEFC";
    attribute INIT_18 of inst : label is "9811000055550000494800005555000009290000292900000909000029290000";
    attribute INIT_19 of inst : label is "FF7F001FFFFF0CFEFFFF303FFFFEE0F00F231F00FCFCFC009185000055550000";
    attribute INIT_1A of inst : label is "0F0F0701FFFFFCF0000200017F7F00FF3F7F1F00FAFEF8005F733F00FC9EFC00";
    attribute INIT_1B of inst : label is "7F723F1FFF1FFEA0FFF97F05FECEFCF87F7F3F05FFFFFE38FFFF7F1CFEFEFCA0";
    attribute INIT_1C of inst : label is "0F1F0000F0F800003F3F0700FCFCE0007F7F1F03FDFEFCC07F271F3AFAFEF8A6";
    attribute INIT_1D of inst : label is "0000000000000000000100000080000003070000C0E00000070F0000E0F00000";
    attribute INIT_1E of inst : label is "3300003F980000F80000003F000000F87F000000FC0000003E13003F3CFC48E0";
    attribute INIT_1F of inst : label is "3F181F00FC38F8003F190300FCC8E000E17E3F3FE070F080FF3E0700E03CFF00";
    attribute INIT_20 of inst : label is "FFC70F3FE0FE013F000000FFFFFFFFFFFFF8FFFFFD83FFFF0000FFFF0000FFFF";
    attribute INIT_21 of inst : label is "FFFFFF0FFFFCFFFFFFFFFFFFFF7F0400FFE00F3FF0FFFFFFFFFFFFF7FFFFFFFF";
    attribute INIT_22 of inst : label is "FFFCF8FF3FFFF0FFFFFF7FFFFC1F7CBE07FF0FC1F0F0FCFFFDE3810CFFE0FFFF";
    attribute INIT_23 of inst : label is "00FF01FFFCFF0FDFFCFF0DFFE0FF3FFF00FFFEFFFFFF7FFFFEFFC30F80FCF03F";
    attribute INIT_24 of inst : label is "FF00FF00FF00FF00FFE0FFFF03FFF8FFFF00FF00007F0000FFF8FFFF00FF00FF";
    attribute INIT_25 of inst : label is "FFFFFF07FFFFFFFF00FFF0FFFF07FFF8FFF0FFFFFFFF0FFFC0FFFFF0FF3FFFFF";
    attribute INIT_26 of inst : label is "F0FF01FF00FF000000000000FF00FF00FFF000FF00FFFFFFFFFFFF00FFF0F8BF";
    attribute INIT_27 of inst : label is "F000FFC0FFFF03FFE080FFFFFFFFFFFFFFFF011FFCC0FFFFFFFFEF0FFF800FFF";
    attribute INIT_28 of inst : label is "00FF00FF00FFFFFF3FFF00FF000FF800FF80FF00FF00FF000000000000C01FFF";
    attribute INIT_29 of inst : label is "00FFFFFF9F0FFFF8FFFFFFFFFFFFFFFFFFFFFFFFF0FFFFF9FFFF000000FF00FF";
    attribute INIT_2A of inst : label is "0000F8FEFFFF010300003F1F000080E0FFFFFFFFFFFFFFFFFFFFFFFFFFFF00FF";
    attribute INIT_2B of inst : label is "C0FCFFFFFFFF0000FCFE0000FFFFFFFF07070000E0F07F1F0000070700C00701";
    attribute INIT_2C of inst : label is "FFFFFFFFFF7FC0FC00F8FEFFFFFF0301F8FE0080E0FFFFFFFFFF000080E03F03";
    attribute INIT_2D of inst : label is "0100FF0F0100FFFFFFFFFFFFFFFFFFFF0F07FF7F1F003F1F0000000000F0F0FF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF00000000FFFFFFFFFFFF7F";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "1F180F00FC0CF8003F301F00F818F0003F1C1900FE1CCC007F383300FC389800";
    attribute INIT_31 of inst : label is "07050000F0D000000F0B0000E0A000001F0A0300FC28E0003F140700F850C000";
    attribute INIT_32 of inst : label is "0003000000C000000003000000C000000303000080E0000001070000C0C00000";
    attribute INIT_33 of inst : label is "0000000000800000000100000000000000010000008000000001000000800000";
    attribute INIT_34 of inst : label is "1F190F00FCFCF8003F331F00F8F8F0003F191C00FEFCFC007F333900FCF8F800";
    attribute INIT_35 of inst : label is "07040000F0F000000F090000E0E000001F0C0300FCF8E0003F190700F8F0C000";
    attribute INIT_36 of inst : label is "070F0700E488F0000F0E03008CC8E0001F1F1900E2C4FC001F110F0086C4F800";
    attribute INIT_37 of inst : label is "03040000E09000000706000090B0000003070300E090E0000704000090900000";
    attribute INIT_38 of inst : label is "7F31001FFE8C00F81F360F00F86CF000FF61007FFF8600FE3F661F00FC66F800";
    attribute INIT_39 of inst : label is "1F070000F8E00000030C0000C03000003F190000FC9800000F140300F028C000";
    attribute INIT_3A of inst : label is "07000000E00000000003000000C000000F000000F00000000005000000E00000";
    attribute INIT_3B of inst : label is "0000000000000000000100000000000000000000000000000003000000800000";
    attribute INIT_3C of inst : label is "6331001FFEFC00F81F390F00F8FCF000E763007FFFFE00FE3F731C00FCFEF800";
    attribute INIT_3D of inst : label is "1B070000F8E00000030D0000C0F00000331F0000FCF800000F190300F0F8C000";
    attribute INIT_3E of inst : label is "3F0F000FFEFC00F80F0E0700F87CF0007F1D003FFFFE00FE1F1C0F00FCFEF800";
    attribute INIT_3F of inst : label is "0F010000F8C0000003060000E0F000001F070000FCF0000007040100F078C000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(5 downto 5),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom6 : if true generate
    attribute INIT_00 of inst : label is "00007FFF00000000E0007F0A0080003FFE260F0100F8000FFFFFFFFF00000000";
    attribute INIT_01 of inst : label is "1EFEF0FFFE1EFFF0FEFEFFFFFEFEFFFF10447EFCFEFF7FFFFE7F7FFE7F7FFFFF";
    attribute INIT_02 of inst : label is "7CF0380100F0001FFC000700004C0006FC000F000098000C00000000387C0000";
    attribute INIT_03 of inst : label is "00000C0030006C0000300000630662436318306360631E06066363701C0C2632";
    attribute INIT_04 of inst : label is "6363736777633030666E03630C0C63633033606030306666333363633663429D";
    attribute INIT_05 of inst : label is "000000000000000000000770330C77776377631C63630C0C6663636E63666360";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "3578DA2F0026007476707B0FC0B40235FEF07B0FC0AC0235FEF07F0FC0FC033F";
    attribute INIT_09 of inst : label is "00000000000000002900050000290041F0007F028080FFFFFF00FF000700007F";
    attribute INIT_0A of inst : label is "FFFF0100000000000000C0E0FF00FFFFFFFF1F030000C0FFFFFF00FF00FF007F";
    attribute INIT_0B of inst : label is "FFFF0001C0F8FFFF1FFFFFFB1FFF00CF00FF00FF00FC00000000C080FFFFFFFF";
    attribute INIT_0C of inst : label is "FFBFF7EF81FF030F0307FEFE3F7FFCFEEFDFE0FF7F7FFFFFDFF7FFFFFDCFFFFF";
    attribute INIT_0D of inst : label is "7F7FF8E0FFFFDFFB7FE7FFFEBF7FF7DFFE3FFFFF3F3F1F3FFEFCBFBFFFFF7FDF";
    attribute INIT_0E of inst : label is "0000F000FF7F0300F8C03F0300000000FFFFF7C77F1FFFFC3F1FFFF00F03FFFE";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "3F1E0F1FFE3CF8807F3C1F01FC78F0F83F1F0F1FFEFCF8807F3F1F01FCF8F0F8";
    attribute INIT_11 of inst : label is "3F1F001FFEFC00FC3F1F7F00FEFCFF001F1F0F00E28CF8001F130303C6CCE090";
    attribute INIT_12 of inst : label is "011F0F00FFFCF000013F1F00FEF8E0C07F301F00FC18F0003F1F0300FEFCE0F8";
    attribute INIT_13 of inst : label is "000000FF000000FFFF0000FFFF0000FF0000F20000004F0000FF7F0000FFFE00";
    attribute INIT_14 of inst : label is "FF3F00FFFFFC00FF7F7F0F07FEFEF0E0F0D0F0F000000000FFFD3F7F80000000";
    attribute INIT_15 of inst : label is "3F1F007FFFFC00FF3F130703FEFEF0E0FE3F00FF7FFC00FF7F790F07FE9EF0E0";
    attribute INIT_16 of inst : label is "F300C0F8F8000000FF0000E0F00000F83C0000FFFE0000FF7F0000FF3C0020FF";
    attribute INIT_17 of inst : label is "FF3F0F07F0F8F0000F1F0F00FFFCF0E0F0F0FFFF1E1EFEFEFFFFFFFFFEFEFEFE";
    attribute INIT_18 of inst : label is "149900005555000049C90000555500007D190000292900000919000029290000";
    attribute INIT_19 of inst : label is "7F3F003FFFFA00FFFF5F007FFEFE00FC07130F00FC0CF8009F930000D5550000";
    attribute INIT_1A of inst : label is "1F090103FFFFF0FC00030000FFFF00FF3E7F070F7EFEE0847F7F1F20FCFEF800";
    attribute INIT_1B of inst : label is "7F7F1F2FFF9FFC7CFFF93F3EFEFEF8F47F7F1F1EFFFFFCBCFFFF3F3DFEFEF878";
    attribute INIT_1C of inst : label is "1F0F0000F8F000003F3F0007FCFC00E07F270F15FEFEF8687F27076DFDFEE052";
    attribute INIT_1D of inst : label is "0000000000000000010000008000000007030000E0C000000F070000F0E00000";
    attribute INIT_1E of inst : label is "3F000038F80000380000001F000000F00F00001CE00000703F01003F7CF80080";
    attribute INIT_1F of inst : label is "3F100F00FC18F0003F19000FFCC800F0C3793F7FE030E0E07F1F030080F2FE00";
    attribute INIT_20 of inst : label is "1FE7001FFFFFF91F3F000000FFFFFF7FFFFCFFFFFFC30000FFFFFFFF0000FFFF";
    attribute INIT_21 of inst : label is "FFFFFF0FFFFFFFFFFFFFFFFFFF3F8300FFF8071FF80FFFFCFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "FFFFFCFF1FFFF8E3FFFF1FFFFE07FF9F1FFF0631FCF8F0FF7EF3000400F8FCFF";
    attribute INIT_23 of inst : label is "00FF007FFFFE07DFCEFC06FFF0FF3F0180FCFFFFFFE1FFE7FCFF0127003FFC1E";
    attribute INIT_24 of inst : label is "FFFFFFFFFF0FFF00FF007FFF00FFFF00FF00FFFF00FF000100C000FF00FF00FF";
    attribute INIT_25 of inst : label is "007FFFF0FFFF00FF00FFFF07FF00FFFFFF00FF00FF0F0000C0FFFFFFFF0FFFFF";
    attribute INIT_26 of inst : label is "FFFF03FF00000000FF00FF00FF00FF00FF00FFC0FFFF00FFFCFFFF00FFFFFEBF";
    attribute INIT_27 of inst : label is "FC00FFE0FFFF013FF880FFFFFFFFFFFF3FFF000FFEF0FFFFFFFFFF0FFFC0FFFF";
    attribute INIT_28 of inst : label is "000000F000FFF0FF0FFF00FF0003FF00FFE0FF00FF00FF000F00000000800F7F";
    attribute INIT_29 of inst : label is "E0FFFFFF9F0FFFFCFFFFFFFFFFFFFFFFFFFFFFFFFCFFFFFFF8FF000000FF000F";
    attribute INIT_2A of inst : label is "3F1F0000033F0000E0E0FFFFFF7F0000FFFFFFFFFFFFFFFFFFFFFFFF3FFF00EF";
    attribute INIT_2B of inst : label is "0000F0FC1F7FF0FCFFFF7F0700C001070000E0F0FFFFFFFF07010000FFFFFFFF";
    attribute INIT_2C of inst : label is "00C0C0FF0000FFFF0000000007070000FFFF0000000080F8010700C0FFFFFFFF";
    attribute INIT_2D of inst : label is "0000FFFFFF3F000000F000FFF0FF07030000FFFFFFFF0000FF3F3F0000000000";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF0F80F800000000FF7F0100";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "1F130300FC34E0003F2C0700F8C8C0003F100F1FFE04F8807F201F01FC08F0F8";
    attribute INIT_31 of inst : label is "07040000F09000000F090000E02000001F0B0000FCE800003F170000F8D00000";
    attribute INIT_32 of inst : label is "03010000C080000003010000C080000003020000E0E0000007050000C0C00000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_34 of inst : label is "1F1F0300FCFCE0003F3F0700F8F8C0003F190F1FFEFCF8807F331F01FCF8F0F8";
    attribute INIT_35 of inst : label is "07070000F0F000000F0F0000E0E000001F0F0000FCF800003F1F0000F8F00000";
    attribute INIT_36 of inst : label is "0F0E0300C498E0000F0E00008CD800001F110F00E28CF8001F1C0303C6CCE090";
    attribute INIT_37 of inst : label is "07060000C8B000000707000098F0000007040000C89000000706000098B00000";
    attribute INIT_38 of inst : label is "7E1F003F7EF800FC3F370300FCECC000FE3F00FF7FFC00FF7F670F07FEE6F0E0";
    attribute INIT_39 of inst : label is "1E00000078000000070B0000E0D000003E07001F7CE000F81F170000F8E80000";
    attribute INIT_3A of inst : label is "07000000E000000000010000008000000F000000F000000003060000C0E00000";
    attribute INIT_3B of inst : label is "0000000000000000000000000000000003000000C00000000003000000800000";
    attribute INIT_3C of inst : label is "631F003FFEF800FC3F3F0300FCFCC000C73100FFFFFC00FF7F730F07FEFEF0E0";
    attribute INIT_3D of inst : label is "19000000F8000000070F0000E0F000003307001FFCE000F81F1F0000F8F80000";
    attribute INIT_3E of inst : label is "1807001FFEF800FC0F0E0100FC7CC000311F007FFFFC00FF3F1C0703FEFEF0E0";
    attribute INIT_3F of inst : label is "0C000000F800000007030000F07000000801000FFCC000F80F070000F8780000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(6 downto 6),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
  rom7 : if true generate
    attribute INIT_00 of inst : label is "00C03EFF00000000C0807F5F0080003FFEFB7F0300F8000FFFFFFFFF00000000";
    attribute INIT_01 of inst : label is "1EFEF0FFFC1E7FF0FEFEFFFFFCFE7FFF00003CFE70FF0EFFFC7F3FFEFFFFAAFF";
    attribute INIT_02 of inst : label is "7CF83E0F00C0000F0CF8060300FC00071CF80C0300F8000F00000000107C0000";
    attribute INIT_03 of inst : label is "003C0C0030306C00003000003E033C4F7F181E637E030E7F3F033E3C0C0C1C63";
    attribute INIT_04 of inst : label is "3E63636F636B3030637C03033F0C63631F637F603F307C631E607E631C7F3CA1";
    attribute INIT_05 of inst : label is "000000000000000000007F38330C633E637F633E63633F0C3C037E7C3E6F7E7E";
    attribute INIT_06 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_07 of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_08 of inst : label is "4A56E875001A00744E786B1D004C0035DEF87B1F005C0035FEF87F1F00FC003F";
    attribute INIT_09 of inst : label is "00000000000000002900050000C6007CF0007F028080FFFFFF00FF0007000000";
    attribute INIT_0A of inst : label is "FFFF0100000000000000C0E0FF81FFFFFFFF3F07000000FE00FF00FF0083007F";
    attribute INIT_0B of inst : label is "FFFF000100F8FFFF07FF7FF900FF008700FF007F000000000000E0C0FFFFC3FF";
    attribute INIT_0C of inst : label is "FFBFF7EFC38F010F0307FCFE7F3FFEFCF7DFF1E3BF7FFFFF9FEFFFFFFEF7FFFF";
    attribute INIT_0D of inst : label is "7F7FFCF0FFFFDFF77F1FFFFFBFBF77EFFFDFFFFF3F3F0F3FFEFEBFBFFFFF7FE1";
    attribute INIT_0E of inst : label is "0000F800FFFF0700FCE03F07F0000F00FFFFFBF77F3FFFFEBF1FFFF81F07FFFE";
    attribute INIT_0F of inst : label is "0000000000000000000000000000000000000000000000000000000000000000";
    attribute INIT_10 of inst : label is "3F1C033FFECCE0FC7F33073FFC38C0FC3F1F033FFEFCE0FC7F3F073FFCF8C0FC";
    attribute INIT_11 of inst : label is "3F1F003FFEFC00FE3F1F3F00FEFCFE001F130307C48CE0F01F13000FC6DC0088";
    attribute INIT_12 of inst : label is "001307037EF8C0F0003F0F037EF080F07F33071FFC98C0D03C1F001F1EFC00FC";
    attribute INIT_13 of inst : label is "0000007F000000FE7F0000FFFE0000FF00007F000000FE001FFE1F00F87FF800";
    attribute INIT_14 of inst : label is "FF1F00FFFFF800FF7F3F031FFEFCC0F8F0F060F000000000FFFD1E7F80800080";
    attribute INIT_15 of inst : label is "3F0F007FFFF800FF3F1F010FFEFCC0F8F81F00FF1FF800FF7F3F031FFEFCC0F8";
    attribute INIT_16 of inst : label is "F3200CF0F00000F8E70030F0F00000781F0200FFFC2000FF3F8008FFF80000FF";
    attribute INIT_17 of inst : label is "FF1F072FF0F8E0C00F1F0703FFF8E0F4F0F07FFF1E1EFCFEFFFF7FFFFEFEFCFE";
    attribute INIT_18 of inst : label is "126600005522000049460000552200004908000029C600000908000029C60000";
    attribute INIT_19 of inst : label is "7F1F007FFFF600FFFF6F00FFFEFC00FE071A030EFC0CF0F89961000055220000";
    attribute INIT_1A of inst : label is "1F090007FFFE00FE03010000FFFE007F383F001F4EFC00E47E7F0F217CFEE0F0";
    attribute INIT_1B of inst : label is "7F7F0755FFFFF07EFEFF0F7E7EFEE0AA7F7F074AFFFFF0BAFFFF0F5DFEFEE052";
    attribute INIT_1C of inst : label is "1F0F0003F8F000C03E1F000F7CF800F07F27032BFFFEE0D47F3F00D7FEFC00EB";
    attribute INIT_1D of inst : label is "010000008000000003000000C000000007000000E00000000F030000F0C00000";
    attribute INIT_1E of inst : label is "1F00003CF000007800000007000000C00300007E800000FC3F00003FE4710008";
    attribute INIT_1F of inst : label is "3F130700FC98C0001C1F001F18F800F8C7790FFCE03080203F1F007F08F3FCC0";
    attribute INIT_20 of inst : label is "FFF71F0700F87F8F00000000FFFFFF3FFFFFFFFFFFE1FFFF0000FFFF0000FFFF";
    attribute INIT_21 of inst : label is "FFFFFFCFFFFFFFFFFFFFFFFFFF1FE301FFFC071FFC00FFFFFFFFFFFFFFFFFFFF";
    attribute INIT_22 of inst : label is "7FFFFEFF0FFFFCE0FFFF0FFFFFC1FF877FC7061B7FFCC0FF3FF8F00FFFFEFFFF";
    attribute INIT_23 of inst : label is "0000C003FFFF876F23E6007FFC1F1F3CC0E0FFFFFF07FF8FFBFF001B000FFFC7";
    attribute INIT_24 of inst : label is "FFFFFFFFFFFFFFFFFFFF1FFF801FFF00FFFFFFFF00FF000F000000FC00FF00FF";
    attribute INIT_25 of inst : label is "000700FF00FF00FFF03FFF00FFF0FFFFFFFFFFFF0F000000F0F8FFFFFF03FFFF";
    attribute INIT_26 of inst : label is "FF000F000000FF00FF00FF00FF00FF00FF00FF00FFF0FFFFE0FFFFF0FFFFFFFF";
    attribute INIT_27 of inst : label is "FF00FFF0FFFF000FFEC0FFFFFFFFFFFF03FF000FFEF8FFFFFFFFFF0FFFF0FFFF";
    attribute INIT_28 of inst : label is "0000000000F800FF03FF00FFF000FF00FFFFFF00FFC0FF03FF00FF000F00033F";
    attribute INIT_29 of inst : label is "FFE0FFFFDF0FFFFEFFFFFFFFFFFFFFFFFFFFFFFFFFFF0FFFC0FF000000000000";
    attribute INIT_2A of inst : label is "0000F0FCFFFF010300003F1F000000C0FFFFFFFFFFFFFFFFFFFFFFFF1FFF8007";
    attribute INIT_2B of inst : label is "00F0FFFFFFFF0000F8FC0000FFFFFFFF07070000C0F0FF3F0000030700800F03";
    attribute INIT_2C of inst : label is "FFFFFFFFFF7F00F000C0F0FFFFFF0301F0FC000000FCFFFFFFFF000000C0FF0F";
    attribute INIT_2D of inst : label is "0300FF7F0F00FFFFFFFFFFFFFFFFFFFF0F07FFFFFF033F1F00000000000000FF";
    attribute INIT_2E of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF000000FF00FFFFFFFFFF";
    attribute INIT_2F of inst : label is "FFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFFF";
    attribute INIT_30 of inst : label is "1F13000FFCB400803F2D0001F8C800F03F13033FFEB4E0FC7F2D073FFCC8C0FC";
    attribute INIT_31 of inst : label is "07070000F0F000000F0F0000E0E000001F0C000FFC9800803F190001F83000F0";
    attribute INIT_32 of inst : label is "03000000C000000003000000C000000003010000E0C0000007030000C0800000";
    attribute INIT_33 of inst : label is "0000000000000000000000000000000001000000800000000100000080000000";
    attribute INIT_34 of inst : label is "1F19000FFCFC00803F330001F8F800F03F1F033FFEFCE0FC7F3F073FFCF8C0FC";
    attribute INIT_35 of inst : label is "07060000F0F000000F0D0000E0E000001F0E000FFC7800803F1C0001F8F000F0";
    attribute INIT_36 of inst : label is "0F0E0000C49800000F090003CCF800901F1C0307C48CE0F01F1C000FC6DC0088";
    attribute INIT_37 of inst : label is "07070000C8F000000703000098E0000007060000C8B000000707000098F00000";
    attribute INIT_38 of inst : label is "6607007F66E000FE3F110007FC8800E0C61F00FF63F800FF7F21031FFE84C0F8";
    attribute INIT_39 of inst : label is "1B00000FD80000F00F050000F0A000003400003F2C0000FC1F090000F8900000";
    attribute INIT_3A of inst : label is "03000000C000000003000000C00000000C000000F000000007030000E0C00000";
    attribute INIT_3B of inst : label is "0100000080000000000000000000000003000000C00000000000000000000000";
    attribute INIT_3C of inst : label is "7F07007FFEE000FE3F190007FCF800E0C71F00FFFFF800FF7F3F031FFEFCC0F8";
    attribute INIT_3D of inst : label is "1F00000FF80000F00F060000F0E000003F00003FFC0000FC1F0C0000F8F00000";
    attribute INIT_3E of inst : label is "1601003F7EE000FE1F0C0001FCF800E0200F007FFFF800FF3F10010FFEFCC0F8";
    attribute INIT_3F of inst : label is "06000007F80000F007020000F06000000E00001FFC0000FC0F060000F8F00000";
  begin
  inst : RAMB16_S1
      --pragma translate_off
      generic map (
        INIT_00 => romgen_str2bv(inst'INIT_00),
        INIT_01 => romgen_str2bv(inst'INIT_01),
        INIT_02 => romgen_str2bv(inst'INIT_02),
        INIT_03 => romgen_str2bv(inst'INIT_03),
        INIT_04 => romgen_str2bv(inst'INIT_04),
        INIT_05 => romgen_str2bv(inst'INIT_05),
        INIT_06 => romgen_str2bv(inst'INIT_06),
        INIT_07 => romgen_str2bv(inst'INIT_07),
        INIT_08 => romgen_str2bv(inst'INIT_08),
        INIT_09 => romgen_str2bv(inst'INIT_09),
        INIT_0A => romgen_str2bv(inst'INIT_0A),
        INIT_0B => romgen_str2bv(inst'INIT_0B),
        INIT_0C => romgen_str2bv(inst'INIT_0C),
        INIT_0D => romgen_str2bv(inst'INIT_0D),
        INIT_0E => romgen_str2bv(inst'INIT_0E),
        INIT_0F => romgen_str2bv(inst'INIT_0F),
        INIT_10 => romgen_str2bv(inst'INIT_10),
        INIT_11 => romgen_str2bv(inst'INIT_11),
        INIT_12 => romgen_str2bv(inst'INIT_12),
        INIT_13 => romgen_str2bv(inst'INIT_13),
        INIT_14 => romgen_str2bv(inst'INIT_14),
        INIT_15 => romgen_str2bv(inst'INIT_15),
        INIT_16 => romgen_str2bv(inst'INIT_16),
        INIT_17 => romgen_str2bv(inst'INIT_17),
        INIT_18 => romgen_str2bv(inst'INIT_18),
        INIT_19 => romgen_str2bv(inst'INIT_19),
        INIT_1A => romgen_str2bv(inst'INIT_1A),
        INIT_1B => romgen_str2bv(inst'INIT_1B),
        INIT_1C => romgen_str2bv(inst'INIT_1C),
        INIT_1D => romgen_str2bv(inst'INIT_1D),
        INIT_1E => romgen_str2bv(inst'INIT_1E),
        INIT_1F => romgen_str2bv(inst'INIT_1F),
        INIT_20 => romgen_str2bv(inst'INIT_20),
        INIT_21 => romgen_str2bv(inst'INIT_21),
        INIT_22 => romgen_str2bv(inst'INIT_22),
        INIT_23 => romgen_str2bv(inst'INIT_23),
        INIT_24 => romgen_str2bv(inst'INIT_24),
        INIT_25 => romgen_str2bv(inst'INIT_25),
        INIT_26 => romgen_str2bv(inst'INIT_26),
        INIT_27 => romgen_str2bv(inst'INIT_27),
        INIT_28 => romgen_str2bv(inst'INIT_28),
        INIT_29 => romgen_str2bv(inst'INIT_29),
        INIT_2A => romgen_str2bv(inst'INIT_2A),
        INIT_2B => romgen_str2bv(inst'INIT_2B),
        INIT_2C => romgen_str2bv(inst'INIT_2C),
        INIT_2D => romgen_str2bv(inst'INIT_2D),
        INIT_2E => romgen_str2bv(inst'INIT_2E),
        INIT_2F => romgen_str2bv(inst'INIT_2F),
        INIT_30 => romgen_str2bv(inst'INIT_30),
        INIT_31 => romgen_str2bv(inst'INIT_31),
        INIT_32 => romgen_str2bv(inst'INIT_32),
        INIT_33 => romgen_str2bv(inst'INIT_33),
        INIT_34 => romgen_str2bv(inst'INIT_34),
        INIT_35 => romgen_str2bv(inst'INIT_35),
        INIT_36 => romgen_str2bv(inst'INIT_36),
        INIT_37 => romgen_str2bv(inst'INIT_37),
        INIT_38 => romgen_str2bv(inst'INIT_38),
        INIT_39 => romgen_str2bv(inst'INIT_39),
        INIT_3A => romgen_str2bv(inst'INIT_3A),
        INIT_3B => romgen_str2bv(inst'INIT_3B),
        INIT_3C => romgen_str2bv(inst'INIT_3C),
        INIT_3D => romgen_str2bv(inst'INIT_3D),
        INIT_3E => romgen_str2bv(inst'INIT_3E),
        INIT_3F => romgen_str2bv(inst'INIT_3F)
        )
      --pragma translate_on
      port map (
        DO   => DATA(7 downto 7),
        ADDR => rom_addr,
        CLK  => CLK,
        DI   => "0",
        EN   => ENA,
        SSR  => '0',
        WE   => '0'
        );
  end generate;
end RTL;
